-------------------------------------------------------
--! @file
--! @brief Translates the Phase from the Phase Accumulator Register to the amplitude of a Sine wave
-------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

--! Receives Phase and returns amplitude of sine wave
entity Sine_LUT is
 port ( address : in std_logic_vector(11 downto 0); --! Phase
    data : out std_logic_vector(11 downto 0)); --! Amplitude
 end entity Sine_LUT;

--! Receives Phase and returns amplitude of sine wave
 architecture arch_Sine_LUT of Sine_LUT is
    type mem is array ( 0 to 2**12 - 1) of std_logic_vector(11 downto 0);
    constant sine_rom : mem := (
    0 => "011111111111",
    1 => "100000000010",
    2 => "100000000101",
    3 => "100000001000",
    4 => "100000001100",
    5 => "100000001111",
    6 => "100000010010",
    7 => "100000010101",
    8 => "100000011000",
    9 => "100000011011",
    10 => "100000011110",
    11 => "100000100010",
    12 => "100000100101",
    13 => "100000101000",
    14 => "100000101011",
    15 => "100000101110",
    16 => "100000110001",
    17 => "100000110100",
    18 => "100000111000",
    19 => "100000111011",
    20 => "100000111110",
    21 => "100001000001",
    22 => "100001000100",
    23 => "100001000111",
    24 => "100001001010",
    25 => "100001001101",
    26 => "100001010001",
    27 => "100001010100",
    28 => "100001010111",
    29 => "100001011010",
    30 => "100001011101",
    31 => "100001100000",
    32 => "100001100011",
    33 => "100001100111",
    34 => "100001101010",
    35 => "100001101101",
    36 => "100001110000",
    37 => "100001110011",
    38 => "100001110110",
    39 => "100001111001",
    40 => "100001111101",
    41 => "100010000000",
    42 => "100010000011",
    43 => "100010000110",
    44 => "100010001001",
    45 => "100010001100",
    46 => "100010001111",
    47 => "100010010010",
    48 => "100010010110",
    49 => "100010011001",
    50 => "100010011100",
    51 => "100010011111",
    52 => "100010100010",
    53 => "100010100101",
    54 => "100010101000",
    55 => "100010101100",
    56 => "100010101111",
    57 => "100010110010",
    58 => "100010110101",
    59 => "100010111000",
    60 => "100010111011",
    61 => "100010111110",
    62 => "100011000001",
    63 => "100011000101",
    64 => "100011001000",
    65 => "100011001011",
    66 => "100011001110",
    67 => "100011010001",
    68 => "100011010100",
    69 => "100011010111",
    70 => "100011011010",
    71 => "100011011110",
    72 => "100011100001",
    73 => "100011100100",
    74 => "100011100111",
    75 => "100011101010",
    76 => "100011101101",
    77 => "100011110000",
    78 => "100011110011",
    79 => "100011110110",
    80 => "100011111010",
    81 => "100011111101",
    82 => "100100000000",
    83 => "100100000011",
    84 => "100100000110",
    85 => "100100001001",
    86 => "100100001100",
    87 => "100100001111",
    88 => "100100010011",
    89 => "100100010110",
    90 => "100100011001",
    91 => "100100011100",
    92 => "100100011111",
    93 => "100100100010",
    94 => "100100100101",
    95 => "100100101000",
    96 => "100100101011",
    97 => "100100101110",
    98 => "100100110010",
    99 => "100100110101",
    100 => "100100111000",
    101 => "100100111011",
    102 => "100100111110",
    103 => "100101000001",
    104 => "100101000100",
    105 => "100101000111",
    106 => "100101001010",
    107 => "100101001110",
    108 => "100101010001",
    109 => "100101010100",
    110 => "100101010111",
    111 => "100101011010",
    112 => "100101011101",
    113 => "100101100000",
    114 => "100101100011",
    115 => "100101100110",
    116 => "100101101001",
    117 => "100101101100",
    118 => "100101110000",
    119 => "100101110011",
    120 => "100101110110",
    121 => "100101111001",
    122 => "100101111100",
    123 => "100101111111",
    124 => "100110000010",
    125 => "100110000101",
    126 => "100110001000",
    127 => "100110001011",
    128 => "100110001110",
    129 => "100110010001",
    130 => "100110010101",
    131 => "100110011000",
    132 => "100110011011",
    133 => "100110011110",
    134 => "100110100001",
    135 => "100110100100",
    136 => "100110100111",
    137 => "100110101010",
    138 => "100110101101",
    139 => "100110110000",
    140 => "100110110011",
    141 => "100110110110",
    142 => "100110111001",
    143 => "100110111100",
    144 => "100111000000",
    145 => "100111000011",
    146 => "100111000110",
    147 => "100111001001",
    148 => "100111001100",
    149 => "100111001111",
    150 => "100111010010",
    151 => "100111010101",
    152 => "100111011000",
    153 => "100111011011",
    154 => "100111011110",
    155 => "100111100001",
    156 => "100111100100",
    157 => "100111100111",
    158 => "100111101010",
    159 => "100111101101",
    160 => "100111110000",
    161 => "100111110011",
    162 => "100111110111",
    163 => "100111111010",
    164 => "100111111101",
    165 => "101000000000",
    166 => "101000000011",
    167 => "101000000110",
    168 => "101000001001",
    169 => "101000001100",
    170 => "101000001111",
    171 => "101000010010",
    172 => "101000010101",
    173 => "101000011000",
    174 => "101000011011",
    175 => "101000011110",
    176 => "101000100001",
    177 => "101000100100",
    178 => "101000100111",
    179 => "101000101010",
    180 => "101000101101",
    181 => "101000110000",
    182 => "101000110011",
    183 => "101000110110",
    184 => "101000111001",
    185 => "101000111100",
    186 => "101000111111",
    187 => "101001000010",
    188 => "101001000101",
    189 => "101001001000",
    190 => "101001001011",
    191 => "101001001110",
    192 => "101001010001",
    193 => "101001010100",
    194 => "101001010111",
    195 => "101001011010",
    196 => "101001011101",
    197 => "101001100000",
    198 => "101001100011",
    199 => "101001100110",
    200 => "101001101001",
    201 => "101001101100",
    202 => "101001101111",
    203 => "101001110010",
    204 => "101001110101",
    205 => "101001111000",
    206 => "101001111011",
    207 => "101001111110",
    208 => "101010000001",
    209 => "101010000100",
    210 => "101010000111",
    211 => "101010001010",
    212 => "101010001101",
    213 => "101010010000",
    214 => "101010010011",
    215 => "101010010110",
    216 => "101010011001",
    217 => "101010011100",
    218 => "101010011111",
    219 => "101010100010",
    220 => "101010100101",
    221 => "101010101000",
    222 => "101010101011",
    223 => "101010101110",
    224 => "101010110001",
    225 => "101010110100",
    226 => "101010110111",
    227 => "101010111010",
    228 => "101010111100",
    229 => "101010111111",
    230 => "101011000010",
    231 => "101011000101",
    232 => "101011001000",
    233 => "101011001011",
    234 => "101011001110",
    235 => "101011010001",
    236 => "101011010100",
    237 => "101011010111",
    238 => "101011011010",
    239 => "101011011101",
    240 => "101011100000",
    241 => "101011100011",
    242 => "101011100110",
    243 => "101011101001",
    244 => "101011101011",
    245 => "101011101110",
    246 => "101011110001",
    247 => "101011110100",
    248 => "101011110111",
    249 => "101011111010",
    250 => "101011111101",
    251 => "101100000000",
    252 => "101100000011",
    253 => "101100000110",
    254 => "101100001001",
    255 => "101100001100",
    256 => "101100001110",
    257 => "101100010001",
    258 => "101100010100",
    259 => "101100010111",
    260 => "101100011010",
    261 => "101100011101",
    262 => "101100100000",
    263 => "101100100011",
    264 => "101100100110",
    265 => "101100101000",
    266 => "101100101011",
    267 => "101100101110",
    268 => "101100110001",
    269 => "101100110100",
    270 => "101100110111",
    271 => "101100111010",
    272 => "101100111101",
    273 => "101100111111",
    274 => "101101000010",
    275 => "101101000101",
    276 => "101101001000",
    277 => "101101001011",
    278 => "101101001110",
    279 => "101101010001",
    280 => "101101010100",
    281 => "101101010110",
    282 => "101101011001",
    283 => "101101011100",
    284 => "101101011111",
    285 => "101101100010",
    286 => "101101100101",
    287 => "101101100111",
    288 => "101101101010",
    289 => "101101101101",
    290 => "101101110000",
    291 => "101101110011",
    292 => "101101110110",
    293 => "101101111000",
    294 => "101101111011",
    295 => "101101111110",
    296 => "101110000001",
    297 => "101110000100",
    298 => "101110000111",
    299 => "101110001001",
    300 => "101110001100",
    301 => "101110001111",
    302 => "101110010010",
    303 => "101110010101",
    304 => "101110010111",
    305 => "101110011010",
    306 => "101110011101",
    307 => "101110100000",
    308 => "101110100011",
    309 => "101110100101",
    310 => "101110101000",
    311 => "101110101011",
    312 => "101110101110",
    313 => "101110110001",
    314 => "101110110011",
    315 => "101110110110",
    316 => "101110111001",
    317 => "101110111100",
    318 => "101110111110",
    319 => "101111000001",
    320 => "101111000100",
    321 => "101111000111",
    322 => "101111001010",
    323 => "101111001100",
    324 => "101111001111",
    325 => "101111010010",
    326 => "101111010101",
    327 => "101111010111",
    328 => "101111011010",
    329 => "101111011101",
    330 => "101111100000",
    331 => "101111100010",
    332 => "101111100101",
    333 => "101111101000",
    334 => "101111101011",
    335 => "101111101101",
    336 => "101111110000",
    337 => "101111110011",
    338 => "101111110110",
    339 => "101111111000",
    340 => "101111111011",
    341 => "101111111110",
    342 => "110000000000",
    343 => "110000000011",
    344 => "110000000110",
    345 => "110000001001",
    346 => "110000001011",
    347 => "110000001110",
    348 => "110000010001",
    349 => "110000010011",
    350 => "110000010110",
    351 => "110000011001",
    352 => "110000011011",
    353 => "110000011110",
    354 => "110000100001",
    355 => "110000100100",
    356 => "110000100110",
    357 => "110000101001",
    358 => "110000101100",
    359 => "110000101110",
    360 => "110000110001",
    361 => "110000110100",
    362 => "110000110110",
    363 => "110000111001",
    364 => "110000111100",
    365 => "110000111110",
    366 => "110001000001",
    367 => "110001000100",
    368 => "110001000110",
    369 => "110001001001",
    370 => "110001001100",
    371 => "110001001110",
    372 => "110001010001",
    373 => "110001010011",
    374 => "110001010110",
    375 => "110001011001",
    376 => "110001011011",
    377 => "110001011110",
    378 => "110001100001",
    379 => "110001100011",
    380 => "110001100110",
    381 => "110001101001",
    382 => "110001101011",
    383 => "110001101110",
    384 => "110001110000",
    385 => "110001110011",
    386 => "110001110110",
    387 => "110001111000",
    388 => "110001111011",
    389 => "110001111101",
    390 => "110010000000",
    391 => "110010000011",
    392 => "110010000101",
    393 => "110010001000",
    394 => "110010001010",
    395 => "110010001101",
    396 => "110010001111",
    397 => "110010010010",
    398 => "110010010101",
    399 => "110010010111",
    400 => "110010011010",
    401 => "110010011100",
    402 => "110010011111",
    403 => "110010100001",
    404 => "110010100100",
    405 => "110010100111",
    406 => "110010101001",
    407 => "110010101100",
    408 => "110010101110",
    409 => "110010110001",
    410 => "110010110011",
    411 => "110010110110",
    412 => "110010111000",
    413 => "110010111011",
    414 => "110010111101",
    415 => "110011000000",
    416 => "110011000011",
    417 => "110011000101",
    418 => "110011001000",
    419 => "110011001010",
    420 => "110011001101",
    421 => "110011001111",
    422 => "110011010010",
    423 => "110011010100",
    424 => "110011010111",
    425 => "110011011001",
    426 => "110011011100",
    427 => "110011011110",
    428 => "110011100001",
    429 => "110011100011",
    430 => "110011100110",
    431 => "110011101000",
    432 => "110011101010",
    433 => "110011101101",
    434 => "110011101111",
    435 => "110011110010",
    436 => "110011110100",
    437 => "110011110111",
    438 => "110011111001",
    439 => "110011111100",
    440 => "110011111110",
    441 => "110100000001",
    442 => "110100000011",
    443 => "110100000110",
    444 => "110100001000",
    445 => "110100001010",
    446 => "110100001101",
    447 => "110100001111",
    448 => "110100010010",
    449 => "110100010100",
    450 => "110100010111",
    451 => "110100011001",
    452 => "110100011011",
    453 => "110100011110",
    454 => "110100100000",
    455 => "110100100011",
    456 => "110100100101",
    457 => "110100100111",
    458 => "110100101010",
    459 => "110100101100",
    460 => "110100101111",
    461 => "110100110001",
    462 => "110100110011",
    463 => "110100110110",
    464 => "110100111000",
    465 => "110100111011",
    466 => "110100111101",
    467 => "110100111111",
    468 => "110101000010",
    469 => "110101000100",
    470 => "110101000110",
    471 => "110101001001",
    472 => "110101001011",
    473 => "110101001101",
    474 => "110101010000",
    475 => "110101010010",
    476 => "110101010100",
    477 => "110101010111",
    478 => "110101011001",
    479 => "110101011011",
    480 => "110101011110",
    481 => "110101100000",
    482 => "110101100010",
    483 => "110101100101",
    484 => "110101100111",
    485 => "110101101001",
    486 => "110101101100",
    487 => "110101101110",
    488 => "110101110000",
    489 => "110101110011",
    490 => "110101110101",
    491 => "110101110111",
    492 => "110101111001",
    493 => "110101111100",
    494 => "110101111110",
    495 => "110110000000",
    496 => "110110000011",
    497 => "110110000101",
    498 => "110110000111",
    499 => "110110001001",
    500 => "110110001100",
    501 => "110110001110",
    502 => "110110010000",
    503 => "110110010010",
    504 => "110110010101",
    505 => "110110010111",
    506 => "110110011001",
    507 => "110110011011",
    508 => "110110011110",
    509 => "110110100000",
    510 => "110110100010",
    511 => "110110100100",
    512 => "110110100111",
    513 => "110110101001",
    514 => "110110101011",
    515 => "110110101101",
    516 => "110110101111",
    517 => "110110110010",
    518 => "110110110100",
    519 => "110110110110",
    520 => "110110111000",
    521 => "110110111010",
    522 => "110110111101",
    523 => "110110111111",
    524 => "110111000001",
    525 => "110111000011",
    526 => "110111000101",
    527 => "110111000111",
    528 => "110111001010",
    529 => "110111001100",
    530 => "110111001110",
    531 => "110111010000",
    532 => "110111010010",
    533 => "110111010100",
    534 => "110111010111",
    535 => "110111011001",
    536 => "110111011011",
    537 => "110111011101",
    538 => "110111011111",
    539 => "110111100001",
    540 => "110111100011",
    541 => "110111100110",
    542 => "110111101000",
    543 => "110111101010",
    544 => "110111101100",
    545 => "110111101110",
    546 => "110111110000",
    547 => "110111110010",
    548 => "110111110100",
    549 => "110111110110",
    550 => "110111111000",
    551 => "110111111011",
    552 => "110111111101",
    553 => "110111111111",
    554 => "111000000001",
    555 => "111000000011",
    556 => "111000000101",
    557 => "111000000111",
    558 => "111000001001",
    559 => "111000001011",
    560 => "111000001101",
    561 => "111000001111",
    562 => "111000010001",
    563 => "111000010011",
    564 => "111000010101",
    565 => "111000010111",
    566 => "111000011001",
    567 => "111000011011",
    568 => "111000011101",
    569 => "111000011111",
    570 => "111000100001",
    571 => "111000100011",
    572 => "111000100101",
    573 => "111000100111",
    574 => "111000101010",
    575 => "111000101011",
    576 => "111000101101",
    577 => "111000101111",
    578 => "111000110001",
    579 => "111000110011",
    580 => "111000110101",
    581 => "111000110111",
    582 => "111000111001",
    583 => "111000111011",
    584 => "111000111101",
    585 => "111000111111",
    586 => "111001000001",
    587 => "111001000011",
    588 => "111001000101",
    589 => "111001000111",
    590 => "111001001001",
    591 => "111001001011",
    592 => "111001001101",
    593 => "111001001111",
    594 => "111001010001",
    595 => "111001010011",
    596 => "111001010101",
    597 => "111001010111",
    598 => "111001011000",
    599 => "111001011010",
    600 => "111001011100",
    601 => "111001011110",
    602 => "111001100000",
    603 => "111001100010",
    604 => "111001100100",
    605 => "111001100110",
    606 => "111001101000",
    607 => "111001101001",
    608 => "111001101011",
    609 => "111001101101",
    610 => "111001101111",
    611 => "111001110001",
    612 => "111001110011",
    613 => "111001110101",
    614 => "111001110110",
    615 => "111001111000",
    616 => "111001111010",
    617 => "111001111100",
    618 => "111001111110",
    619 => "111010000000",
    620 => "111010000001",
    621 => "111010000011",
    622 => "111010000101",
    623 => "111010000111",
    624 => "111010001001",
    625 => "111010001011",
    626 => "111010001100",
    627 => "111010001110",
    628 => "111010010000",
    629 => "111010010010",
    630 => "111010010100",
    631 => "111010010101",
    632 => "111010010111",
    633 => "111010011001",
    634 => "111010011011",
    635 => "111010011100",
    636 => "111010011110",
    637 => "111010100000",
    638 => "111010100010",
    639 => "111010100011",
    640 => "111010100101",
    641 => "111010100111",
    642 => "111010101001",
    643 => "111010101010",
    644 => "111010101100",
    645 => "111010101110",
    646 => "111010110000",
    647 => "111010110001",
    648 => "111010110011",
    649 => "111010110101",
    650 => "111010110110",
    651 => "111010111000",
    652 => "111010111010",
    653 => "111010111100",
    654 => "111010111101",
    655 => "111010111111",
    656 => "111011000001",
    657 => "111011000010",
    658 => "111011000100",
    659 => "111011000110",
    660 => "111011000111",
    661 => "111011001001",
    662 => "111011001011",
    663 => "111011001100",
    664 => "111011001110",
    665 => "111011010000",
    666 => "111011010001",
    667 => "111011010011",
    668 => "111011010100",
    669 => "111011010110",
    670 => "111011011000",
    671 => "111011011001",
    672 => "111011011011",
    673 => "111011011101",
    674 => "111011011110",
    675 => "111011100000",
    676 => "111011100001",
    677 => "111011100011",
    678 => "111011100101",
    679 => "111011100110",
    680 => "111011101000",
    681 => "111011101001",
    682 => "111011101011",
    683 => "111011101100",
    684 => "111011101110",
    685 => "111011110000",
    686 => "111011110001",
    687 => "111011110011",
    688 => "111011110100",
    689 => "111011110110",
    690 => "111011110111",
    691 => "111011111001",
    692 => "111011111010",
    693 => "111011111100",
    694 => "111011111101",
    695 => "111011111111",
    696 => "111100000000",
    697 => "111100000010",
    698 => "111100000011",
    699 => "111100000101",
    700 => "111100000110",
    701 => "111100001000",
    702 => "111100001001",
    703 => "111100001011",
    704 => "111100001100",
    705 => "111100001110",
    706 => "111100001111",
    707 => "111100010001",
    708 => "111100010010",
    709 => "111100010100",
    710 => "111100010101",
    711 => "111100010111",
    712 => "111100011000",
    713 => "111100011010",
    714 => "111100011011",
    715 => "111100011100",
    716 => "111100011110",
    717 => "111100011111",
    718 => "111100100001",
    719 => "111100100010",
    720 => "111100100100",
    721 => "111100100101",
    722 => "111100100110",
    723 => "111100101000",
    724 => "111100101001",
    725 => "111100101011",
    726 => "111100101100",
    727 => "111100101101",
    728 => "111100101111",
    729 => "111100110000",
    730 => "111100110001",
    731 => "111100110011",
    732 => "111100110100",
    733 => "111100110110",
    734 => "111100110111",
    735 => "111100111000",
    736 => "111100111010",
    737 => "111100111011",
    738 => "111100111100",
    739 => "111100111110",
    740 => "111100111111",
    741 => "111101000000",
    742 => "111101000010",
    743 => "111101000011",
    744 => "111101000100",
    745 => "111101000110",
    746 => "111101000111",
    747 => "111101001000",
    748 => "111101001001",
    749 => "111101001011",
    750 => "111101001100",
    751 => "111101001101",
    752 => "111101001111",
    753 => "111101010000",
    754 => "111101010001",
    755 => "111101010010",
    756 => "111101010100",
    757 => "111101010101",
    758 => "111101010110",
    759 => "111101010111",
    760 => "111101011001",
    761 => "111101011010",
    762 => "111101011011",
    763 => "111101011100",
    764 => "111101011110",
    765 => "111101011111",
    766 => "111101100000",
    767 => "111101100001",
    768 => "111101100010",
    769 => "111101100100",
    770 => "111101100101",
    771 => "111101100110",
    772 => "111101100111",
    773 => "111101101000",
    774 => "111101101001",
    775 => "111101101011",
    776 => "111101101100",
    777 => "111101101101",
    778 => "111101101110",
    779 => "111101101111",
    780 => "111101110000",
    781 => "111101110010",
    782 => "111101110011",
    783 => "111101110100",
    784 => "111101110101",
    785 => "111101110110",
    786 => "111101110111",
    787 => "111101111000",
    788 => "111101111001",
    789 => "111101111011",
    790 => "111101111100",
    791 => "111101111101",
    792 => "111101111110",
    793 => "111101111111",
    794 => "111110000000",
    795 => "111110000001",
    796 => "111110000010",
    797 => "111110000011",
    798 => "111110000100",
    799 => "111110000101",
    800 => "111110000111",
    801 => "111110001000",
    802 => "111110001001",
    803 => "111110001010",
    804 => "111110001011",
    805 => "111110001100",
    806 => "111110001101",
    807 => "111110001110",
    808 => "111110001111",
    809 => "111110010000",
    810 => "111110010001",
    811 => "111110010010",
    812 => "111110010011",
    813 => "111110010100",
    814 => "111110010101",
    815 => "111110010110",
    816 => "111110010111",
    817 => "111110011000",
    818 => "111110011001",
    819 => "111110011010",
    820 => "111110011011",
    821 => "111110011100",
    822 => "111110011101",
    823 => "111110011110",
    824 => "111110011111",
    825 => "111110100000",
    826 => "111110100000",
    827 => "111110100001",
    828 => "111110100010",
    829 => "111110100011",
    830 => "111110100100",
    831 => "111110100101",
    832 => "111110100110",
    833 => "111110100111",
    834 => "111110101000",
    835 => "111110101001",
    836 => "111110101010",
    837 => "111110101011",
    838 => "111110101011",
    839 => "111110101100",
    840 => "111110101101",
    841 => "111110101110",
    842 => "111110101111",
    843 => "111110110000",
    844 => "111110110001",
    845 => "111110110001",
    846 => "111110110010",
    847 => "111110110011",
    848 => "111110110100",
    849 => "111110110101",
    850 => "111110110110",
    851 => "111110110111",
    852 => "111110110111",
    853 => "111110111000",
    854 => "111110111001",
    855 => "111110111010",
    856 => "111110111011",
    857 => "111110111011",
    858 => "111110111100",
    859 => "111110111101",
    860 => "111110111110",
    861 => "111110111111",
    862 => "111110111111",
    863 => "111111000000",
    864 => "111111000001",
    865 => "111111000010",
    866 => "111111000010",
    867 => "111111000011",
    868 => "111111000100",
    869 => "111111000101",
    870 => "111111000101",
    871 => "111111000110",
    872 => "111111000111",
    873 => "111111001000",
    874 => "111111001000",
    875 => "111111001001",
    876 => "111111001010",
    877 => "111111001010",
    878 => "111111001011",
    879 => "111111001100",
    880 => "111111001100",
    881 => "111111001101",
    882 => "111111001110",
    883 => "111111001110",
    884 => "111111001111",
    885 => "111111010000",
    886 => "111111010000",
    887 => "111111010001",
    888 => "111111010010",
    889 => "111111010010",
    890 => "111111010011",
    891 => "111111010100",
    892 => "111111010100",
    893 => "111111010101",
    894 => "111111010110",
    895 => "111111010110",
    896 => "111111010111",
    897 => "111111010111",
    898 => "111111011000",
    899 => "111111011001",
    900 => "111111011001",
    901 => "111111011010",
    902 => "111111011010",
    903 => "111111011011",
    904 => "111111011100",
    905 => "111111011100",
    906 => "111111011101",
    907 => "111111011101",
    908 => "111111011110",
    909 => "111111011110",
    910 => "111111011111",
    911 => "111111100000",
    912 => "111111100000",
    913 => "111111100001",
    914 => "111111100001",
    915 => "111111100010",
    916 => "111111100010",
    917 => "111111100011",
    918 => "111111100011",
    919 => "111111100100",
    920 => "111111100100",
    921 => "111111100101",
    922 => "111111100101",
    923 => "111111100110",
    924 => "111111100110",
    925 => "111111100111",
    926 => "111111100111",
    927 => "111111101000",
    928 => "111111101000",
    929 => "111111101000",
    930 => "111111101001",
    931 => "111111101001",
    932 => "111111101010",
    933 => "111111101010",
    934 => "111111101011",
    935 => "111111101011",
    936 => "111111101100",
    937 => "111111101100",
    938 => "111111101100",
    939 => "111111101101",
    940 => "111111101101",
    941 => "111111101110",
    942 => "111111101110",
    943 => "111111101110",
    944 => "111111101111",
    945 => "111111101111",
    946 => "111111110000",
    947 => "111111110000",
    948 => "111111110000",
    949 => "111111110001",
    950 => "111111110001",
    951 => "111111110001",
    952 => "111111110010",
    953 => "111111110010",
    954 => "111111110010",
    955 => "111111110011",
    956 => "111111110011",
    957 => "111111110011",
    958 => "111111110100",
    959 => "111111110100",
    960 => "111111110100",
    961 => "111111110101",
    962 => "111111110101",
    963 => "111111110101",
    964 => "111111110110",
    965 => "111111110110",
    966 => "111111110110",
    967 => "111111110110",
    968 => "111111110111",
    969 => "111111110111",
    970 => "111111110111",
    971 => "111111110111",
    972 => "111111111000",
    973 => "111111111000",
    974 => "111111111000",
    975 => "111111111000",
    976 => "111111111001",
    977 => "111111111001",
    978 => "111111111001",
    979 => "111111111001",
    980 => "111111111010",
    981 => "111111111010",
    982 => "111111111010",
    983 => "111111111010",
    984 => "111111111010",
    985 => "111111111011",
    986 => "111111111011",
    987 => "111111111011",
    988 => "111111111011",
    989 => "111111111011",
    990 => "111111111011",
    991 => "111111111100",
    992 => "111111111100",
    993 => "111111111100",
    994 => "111111111100",
    995 => "111111111100",
    996 => "111111111100",
    997 => "111111111100",
    998 => "111111111101",
    999 => "111111111101",
    1000 => "111111111101",
    1001 => "111111111101",
    1002 => "111111111101",
    1003 => "111111111101",
    1004 => "111111111101",
    1005 => "111111111101",
    1006 => "111111111101",
    1007 => "111111111101",
    1008 => "111111111110",
    1009 => "111111111110",
    1010 => "111111111110",
    1011 => "111111111110",
    1012 => "111111111110",
    1013 => "111111111110",
    1014 => "111111111110",
    1015 => "111111111110",
    1016 => "111111111110",
    1017 => "111111111110",
    1018 => "111111111110",
    1019 => "111111111110",
    1020 => "111111111110",
    1021 => "111111111110",
    1022 => "111111111110",
    1023 => "111111111110",
    1024 => "111111111110",
    1025 => "111111111110",
    1026 => "111111111110",
    1027 => "111111111110",
    1028 => "111111111110",
    1029 => "111111111110",
    1030 => "111111111110",
    1031 => "111111111110",
    1032 => "111111111110",
    1033 => "111111111110",
    1034 => "111111111110",
    1035 => "111111111110",
    1036 => "111111111110",
    1037 => "111111111110",
    1038 => "111111111110",
    1039 => "111111111110",
    1040 => "111111111110",
    1041 => "111111111101",
    1042 => "111111111101",
    1043 => "111111111101",
    1044 => "111111111101",
    1045 => "111111111101",
    1046 => "111111111101",
    1047 => "111111111101",
    1048 => "111111111101",
    1049 => "111111111101",
    1050 => "111111111101",
    1051 => "111111111100",
    1052 => "111111111100",
    1053 => "111111111100",
    1054 => "111111111100",
    1055 => "111111111100",
    1056 => "111111111100",
    1057 => "111111111100",
    1058 => "111111111011",
    1059 => "111111111011",
    1060 => "111111111011",
    1061 => "111111111011",
    1062 => "111111111011",
    1063 => "111111111011",
    1064 => "111111111010",
    1065 => "111111111010",
    1066 => "111111111010",
    1067 => "111111111010",
    1068 => "111111111010",
    1069 => "111111111001",
    1070 => "111111111001",
    1071 => "111111111001",
    1072 => "111111111001",
    1073 => "111111111000",
    1074 => "111111111000",
    1075 => "111111111000",
    1076 => "111111111000",
    1077 => "111111110111",
    1078 => "111111110111",
    1079 => "111111110111",
    1080 => "111111110111",
    1081 => "111111110110",
    1082 => "111111110110",
    1083 => "111111110110",
    1084 => "111111110110",
    1085 => "111111110101",
    1086 => "111111110101",
    1087 => "111111110101",
    1088 => "111111110100",
    1089 => "111111110100",
    1090 => "111111110100",
    1091 => "111111110011",
    1092 => "111111110011",
    1093 => "111111110011",
    1094 => "111111110010",
    1095 => "111111110010",
    1096 => "111111110010",
    1097 => "111111110001",
    1098 => "111111110001",
    1099 => "111111110001",
    1100 => "111111110000",
    1101 => "111111110000",
    1102 => "111111110000",
    1103 => "111111101111",
    1104 => "111111101111",
    1105 => "111111101110",
    1106 => "111111101110",
    1107 => "111111101110",
    1108 => "111111101101",
    1109 => "111111101101",
    1110 => "111111101100",
    1111 => "111111101100",
    1112 => "111111101100",
    1113 => "111111101011",
    1114 => "111111101011",
    1115 => "111111101010",
    1116 => "111111101010",
    1117 => "111111101001",
    1118 => "111111101001",
    1119 => "111111101000",
    1120 => "111111101000",
    1121 => "111111101000",
    1122 => "111111100111",
    1123 => "111111100111",
    1124 => "111111100110",
    1125 => "111111100110",
    1126 => "111111100101",
    1127 => "111111100101",
    1128 => "111111100100",
    1129 => "111111100100",
    1130 => "111111100011",
    1131 => "111111100011",
    1132 => "111111100010",
    1133 => "111111100010",
    1134 => "111111100001",
    1135 => "111111100001",
    1136 => "111111100000",
    1137 => "111111100000",
    1138 => "111111011111",
    1139 => "111111011110",
    1140 => "111111011110",
    1141 => "111111011101",
    1142 => "111111011101",
    1143 => "111111011100",
    1144 => "111111011100",
    1145 => "111111011011",
    1146 => "111111011010",
    1147 => "111111011010",
    1148 => "111111011001",
    1149 => "111111011001",
    1150 => "111111011000",
    1151 => "111111010111",
    1152 => "111111010111",
    1153 => "111111010110",
    1154 => "111111010110",
    1155 => "111111010101",
    1156 => "111111010100",
    1157 => "111111010100",
    1158 => "111111010011",
    1159 => "111111010010",
    1160 => "111111010010",
    1161 => "111111010001",
    1162 => "111111010000",
    1163 => "111111010000",
    1164 => "111111001111",
    1165 => "111111001110",
    1166 => "111111001110",
    1167 => "111111001101",
    1168 => "111111001100",
    1169 => "111111001100",
    1170 => "111111001011",
    1171 => "111111001010",
    1172 => "111111001010",
    1173 => "111111001001",
    1174 => "111111001000",
    1175 => "111111001000",
    1176 => "111111000111",
    1177 => "111111000110",
    1178 => "111111000101",
    1179 => "111111000101",
    1180 => "111111000100",
    1181 => "111111000011",
    1182 => "111111000010",
    1183 => "111111000010",
    1184 => "111111000001",
    1185 => "111111000000",
    1186 => "111110111111",
    1187 => "111110111111",
    1188 => "111110111110",
    1189 => "111110111101",
    1190 => "111110111100",
    1191 => "111110111011",
    1192 => "111110111011",
    1193 => "111110111010",
    1194 => "111110111001",
    1195 => "111110111000",
    1196 => "111110110111",
    1197 => "111110110111",
    1198 => "111110110110",
    1199 => "111110110101",
    1200 => "111110110100",
    1201 => "111110110011",
    1202 => "111110110010",
    1203 => "111110110001",
    1204 => "111110110001",
    1205 => "111110110000",
    1206 => "111110101111",
    1207 => "111110101110",
    1208 => "111110101101",
    1209 => "111110101100",
    1210 => "111110101011",
    1211 => "111110101011",
    1212 => "111110101010",
    1213 => "111110101001",
    1214 => "111110101000",
    1215 => "111110100111",
    1216 => "111110100110",
    1217 => "111110100101",
    1218 => "111110100100",
    1219 => "111110100011",
    1220 => "111110100010",
    1221 => "111110100001",
    1222 => "111110100000",
    1223 => "111110100000",
    1224 => "111110011111",
    1225 => "111110011110",
    1226 => "111110011101",
    1227 => "111110011100",
    1228 => "111110011011",
    1229 => "111110011010",
    1230 => "111110011001",
    1231 => "111110011000",
    1232 => "111110010111",
    1233 => "111110010110",
    1234 => "111110010101",
    1235 => "111110010100",
    1236 => "111110010011",
    1237 => "111110010010",
    1238 => "111110010001",
    1239 => "111110010000",
    1240 => "111110001111",
    1241 => "111110001110",
    1242 => "111110001101",
    1243 => "111110001100",
    1244 => "111110001011",
    1245 => "111110001010",
    1246 => "111110001001",
    1247 => "111110001000",
    1248 => "111110000111",
    1249 => "111110000101",
    1250 => "111110000100",
    1251 => "111110000011",
    1252 => "111110000010",
    1253 => "111110000001",
    1254 => "111110000000",
    1255 => "111101111111",
    1256 => "111101111110",
    1257 => "111101111101",
    1258 => "111101111100",
    1259 => "111101111011",
    1260 => "111101111001",
    1261 => "111101111000",
    1262 => "111101110111",
    1263 => "111101110110",
    1264 => "111101110101",
    1265 => "111101110100",
    1266 => "111101110011",
    1267 => "111101110010",
    1268 => "111101110000",
    1269 => "111101101111",
    1270 => "111101101110",
    1271 => "111101101101",
    1272 => "111101101100",
    1273 => "111101101011",
    1274 => "111101101001",
    1275 => "111101101000",
    1276 => "111101100111",
    1277 => "111101100110",
    1278 => "111101100101",
    1279 => "111101100100",
    1280 => "111101100010",
    1281 => "111101100001",
    1282 => "111101100000",
    1283 => "111101011111",
    1284 => "111101011110",
    1285 => "111101011100",
    1286 => "111101011011",
    1287 => "111101011010",
    1288 => "111101011001",
    1289 => "111101010111",
    1290 => "111101010110",
    1291 => "111101010101",
    1292 => "111101010100",
    1293 => "111101010010",
    1294 => "111101010001",
    1295 => "111101010000",
    1296 => "111101001111",
    1297 => "111101001101",
    1298 => "111101001100",
    1299 => "111101001011",
    1300 => "111101001001",
    1301 => "111101001000",
    1302 => "111101000111",
    1303 => "111101000110",
    1304 => "111101000100",
    1305 => "111101000011",
    1306 => "111101000010",
    1307 => "111101000000",
    1308 => "111100111111",
    1309 => "111100111110",
    1310 => "111100111100",
    1311 => "111100111011",
    1312 => "111100111010",
    1313 => "111100111000",
    1314 => "111100110111",
    1315 => "111100110110",
    1316 => "111100110100",
    1317 => "111100110011",
    1318 => "111100110001",
    1319 => "111100110000",
    1320 => "111100101111",
    1321 => "111100101101",
    1322 => "111100101100",
    1323 => "111100101011",
    1324 => "111100101001",
    1325 => "111100101000",
    1326 => "111100100110",
    1327 => "111100100101",
    1328 => "111100100100",
    1329 => "111100100010",
    1330 => "111100100001",
    1331 => "111100011111",
    1332 => "111100011110",
    1333 => "111100011100",
    1334 => "111100011011",
    1335 => "111100011010",
    1336 => "111100011000",
    1337 => "111100010111",
    1338 => "111100010101",
    1339 => "111100010100",
    1340 => "111100010010",
    1341 => "111100010001",
    1342 => "111100001111",
    1343 => "111100001110",
    1344 => "111100001100",
    1345 => "111100001011",
    1346 => "111100001001",
    1347 => "111100001000",
    1348 => "111100000110",
    1349 => "111100000101",
    1350 => "111100000011",
    1351 => "111100000010",
    1352 => "111100000000",
    1353 => "111011111111",
    1354 => "111011111101",
    1355 => "111011111100",
    1356 => "111011111010",
    1357 => "111011111001",
    1358 => "111011110111",
    1359 => "111011110110",
    1360 => "111011110100",
    1361 => "111011110011",
    1362 => "111011110001",
    1363 => "111011110000",
    1364 => "111011101110",
    1365 => "111011101100",
    1366 => "111011101011",
    1367 => "111011101001",
    1368 => "111011101000",
    1369 => "111011100110",
    1370 => "111011100101",
    1371 => "111011100011",
    1372 => "111011100001",
    1373 => "111011100000",
    1374 => "111011011110",
    1375 => "111011011101",
    1376 => "111011011011",
    1377 => "111011011001",
    1378 => "111011011000",
    1379 => "111011010110",
    1380 => "111011010100",
    1381 => "111011010011",
    1382 => "111011010001",
    1383 => "111011010000",
    1384 => "111011001110",
    1385 => "111011001100",
    1386 => "111011001011",
    1387 => "111011001001",
    1388 => "111011000111",
    1389 => "111011000110",
    1390 => "111011000100",
    1391 => "111011000010",
    1392 => "111011000001",
    1393 => "111010111111",
    1394 => "111010111101",
    1395 => "111010111100",
    1396 => "111010111010",
    1397 => "111010111000",
    1398 => "111010110110",
    1399 => "111010110101",
    1400 => "111010110011",
    1401 => "111010110001",
    1402 => "111010110000",
    1403 => "111010101110",
    1404 => "111010101100",
    1405 => "111010101010",
    1406 => "111010101001",
    1407 => "111010100111",
    1408 => "111010100101",
    1409 => "111010100011",
    1410 => "111010100010",
    1411 => "111010100000",
    1412 => "111010011110",
    1413 => "111010011100",
    1414 => "111010011011",
    1415 => "111010011001",
    1416 => "111010010111",
    1417 => "111010010101",
    1418 => "111010010100",
    1419 => "111010010010",
    1420 => "111010010000",
    1421 => "111010001110",
    1422 => "111010001100",
    1423 => "111010001011",
    1424 => "111010001001",
    1425 => "111010000111",
    1426 => "111010000101",
    1427 => "111010000011",
    1428 => "111010000001",
    1429 => "111010000000",
    1430 => "111001111110",
    1431 => "111001111100",
    1432 => "111001111010",
    1433 => "111001111000",
    1434 => "111001110110",
    1435 => "111001110101",
    1436 => "111001110011",
    1437 => "111001110001",
    1438 => "111001101111",
    1439 => "111001101101",
    1440 => "111001101011",
    1441 => "111001101001",
    1442 => "111001101000",
    1443 => "111001100110",
    1444 => "111001100100",
    1445 => "111001100010",
    1446 => "111001100000",
    1447 => "111001011110",
    1448 => "111001011100",
    1449 => "111001011010",
    1450 => "111001011000",
    1451 => "111001010111",
    1452 => "111001010101",
    1453 => "111001010011",
    1454 => "111001010001",
    1455 => "111001001111",
    1456 => "111001001101",
    1457 => "111001001011",
    1458 => "111001001001",
    1459 => "111001000111",
    1460 => "111001000101",
    1461 => "111001000011",
    1462 => "111001000001",
    1463 => "111000111111",
    1464 => "111000111101",
    1465 => "111000111011",
    1466 => "111000111001",
    1467 => "111000110111",
    1468 => "111000110101",
    1469 => "111000110011",
    1470 => "111000110001",
    1471 => "111000101111",
    1472 => "111000101101",
    1473 => "111000101011",
    1474 => "111000101010",
    1475 => "111000100111",
    1476 => "111000100101",
    1477 => "111000100011",
    1478 => "111000100001",
    1479 => "111000011111",
    1480 => "111000011101",
    1481 => "111000011011",
    1482 => "111000011001",
    1483 => "111000010111",
    1484 => "111000010101",
    1485 => "111000010011",
    1486 => "111000010001",
    1487 => "111000001111",
    1488 => "111000001101",
    1489 => "111000001011",
    1490 => "111000001001",
    1491 => "111000000111",
    1492 => "111000000101",
    1493 => "111000000011",
    1494 => "111000000001",
    1495 => "110111111111",
    1496 => "110111111101",
    1497 => "110111111011",
    1498 => "110111111000",
    1499 => "110111110110",
    1500 => "110111110100",
    1501 => "110111110010",
    1502 => "110111110000",
    1503 => "110111101110",
    1504 => "110111101100",
    1505 => "110111101010",
    1506 => "110111101000",
    1507 => "110111100110",
    1508 => "110111100011",
    1509 => "110111100001",
    1510 => "110111011111",
    1511 => "110111011101",
    1512 => "110111011011",
    1513 => "110111011001",
    1514 => "110111010111",
    1515 => "110111010100",
    1516 => "110111010010",
    1517 => "110111010000",
    1518 => "110111001110",
    1519 => "110111001100",
    1520 => "110111001010",
    1521 => "110111000111",
    1522 => "110111000101",
    1523 => "110111000011",
    1524 => "110111000001",
    1525 => "110110111111",
    1526 => "110110111101",
    1527 => "110110111010",
    1528 => "110110111000",
    1529 => "110110110110",
    1530 => "110110110100",
    1531 => "110110110010",
    1532 => "110110101111",
    1533 => "110110101101",
    1534 => "110110101011",
    1535 => "110110101001",
    1536 => "110110100111",
    1537 => "110110100100",
    1538 => "110110100010",
    1539 => "110110100000",
    1540 => "110110011110",
    1541 => "110110011011",
    1542 => "110110011001",
    1543 => "110110010111",
    1544 => "110110010101",
    1545 => "110110010010",
    1546 => "110110010000",
    1547 => "110110001110",
    1548 => "110110001100",
    1549 => "110110001001",
    1550 => "110110000111",
    1551 => "110110000101",
    1552 => "110110000011",
    1553 => "110110000000",
    1554 => "110101111110",
    1555 => "110101111100",
    1556 => "110101111001",
    1557 => "110101110111",
    1558 => "110101110101",
    1559 => "110101110011",
    1560 => "110101110000",
    1561 => "110101101110",
    1562 => "110101101100",
    1563 => "110101101001",
    1564 => "110101100111",
    1565 => "110101100101",
    1566 => "110101100010",
    1567 => "110101100000",
    1568 => "110101011110",
    1569 => "110101011011",
    1570 => "110101011001",
    1571 => "110101010111",
    1572 => "110101010100",
    1573 => "110101010010",
    1574 => "110101010000",
    1575 => "110101001101",
    1576 => "110101001011",
    1577 => "110101001001",
    1578 => "110101000110",
    1579 => "110101000100",
    1580 => "110101000010",
    1581 => "110100111111",
    1582 => "110100111101",
    1583 => "110100111011",
    1584 => "110100111000",
    1585 => "110100110110",
    1586 => "110100110011",
    1587 => "110100110001",
    1588 => "110100101111",
    1589 => "110100101100",
    1590 => "110100101010",
    1591 => "110100100111",
    1592 => "110100100101",
    1593 => "110100100011",
    1594 => "110100100000",
    1595 => "110100011110",
    1596 => "110100011011",
    1597 => "110100011001",
    1598 => "110100010111",
    1599 => "110100010100",
    1600 => "110100010010",
    1601 => "110100001111",
    1602 => "110100001101",
    1603 => "110100001010",
    1604 => "110100001000",
    1605 => "110100000110",
    1606 => "110100000011",
    1607 => "110100000001",
    1608 => "110011111110",
    1609 => "110011111100",
    1610 => "110011111001",
    1611 => "110011110111",
    1612 => "110011110100",
    1613 => "110011110010",
    1614 => "110011101111",
    1615 => "110011101101",
    1616 => "110011101010",
    1617 => "110011101000",
    1618 => "110011100110",
    1619 => "110011100011",
    1620 => "110011100001",
    1621 => "110011011110",
    1622 => "110011011100",
    1623 => "110011011001",
    1624 => "110011010111",
    1625 => "110011010100",
    1626 => "110011010010",
    1627 => "110011001111",
    1628 => "110011001101",
    1629 => "110011001010",
    1630 => "110011001000",
    1631 => "110011000101",
    1632 => "110011000011",
    1633 => "110011000000",
    1634 => "110010111101",
    1635 => "110010111011",
    1636 => "110010111000",
    1637 => "110010110110",
    1638 => "110010110011",
    1639 => "110010110001",
    1640 => "110010101110",
    1641 => "110010101100",
    1642 => "110010101001",
    1643 => "110010100111",
    1644 => "110010100100",
    1645 => "110010100001",
    1646 => "110010011111",
    1647 => "110010011100",
    1648 => "110010011010",
    1649 => "110010010111",
    1650 => "110010010101",
    1651 => "110010010010",
    1652 => "110010001111",
    1653 => "110010001101",
    1654 => "110010001010",
    1655 => "110010001000",
    1656 => "110010000101",
    1657 => "110010000011",
    1658 => "110010000000",
    1659 => "110001111101",
    1660 => "110001111011",
    1661 => "110001111000",
    1662 => "110001110110",
    1663 => "110001110011",
    1664 => "110001110000",
    1665 => "110001101110",
    1666 => "110001101011",
    1667 => "110001101001",
    1668 => "110001100110",
    1669 => "110001100011",
    1670 => "110001100001",
    1671 => "110001011110",
    1672 => "110001011011",
    1673 => "110001011001",
    1674 => "110001010110",
    1675 => "110001010011",
    1676 => "110001010001",
    1677 => "110001001110",
    1678 => "110001001100",
    1679 => "110001001001",
    1680 => "110001000110",
    1681 => "110001000100",
    1682 => "110001000001",
    1683 => "110000111110",
    1684 => "110000111100",
    1685 => "110000111001",
    1686 => "110000110110",
    1687 => "110000110100",
    1688 => "110000110001",
    1689 => "110000101110",
    1690 => "110000101100",
    1691 => "110000101001",
    1692 => "110000100110",
    1693 => "110000100100",
    1694 => "110000100001",
    1695 => "110000011110",
    1696 => "110000011011",
    1697 => "110000011001",
    1698 => "110000010110",
    1699 => "110000010011",
    1700 => "110000010001",
    1701 => "110000001110",
    1702 => "110000001011",
    1703 => "110000001001",
    1704 => "110000000110",
    1705 => "110000000011",
    1706 => "110000000000",
    1707 => "101111111110",
    1708 => "101111111011",
    1709 => "101111111000",
    1710 => "101111110110",
    1711 => "101111110011",
    1712 => "101111110000",
    1713 => "101111101101",
    1714 => "101111101011",
    1715 => "101111101000",
    1716 => "101111100101",
    1717 => "101111100010",
    1718 => "101111100000",
    1719 => "101111011101",
    1720 => "101111011010",
    1721 => "101111010111",
    1722 => "101111010101",
    1723 => "101111010010",
    1724 => "101111001111",
    1725 => "101111001100",
    1726 => "101111001010",
    1727 => "101111000111",
    1728 => "101111000100",
    1729 => "101111000001",
    1730 => "101110111110",
    1731 => "101110111100",
    1732 => "101110111001",
    1733 => "101110110110",
    1734 => "101110110011",
    1735 => "101110110001",
    1736 => "101110101110",
    1737 => "101110101011",
    1738 => "101110101000",
    1739 => "101110100101",
    1740 => "101110100011",
    1741 => "101110100000",
    1742 => "101110011101",
    1743 => "101110011010",
    1744 => "101110010111",
    1745 => "101110010101",
    1746 => "101110010010",
    1747 => "101110001111",
    1748 => "101110001100",
    1749 => "101110001001",
    1750 => "101110000111",
    1751 => "101110000100",
    1752 => "101110000001",
    1753 => "101101111110",
    1754 => "101101111011",
    1755 => "101101111000",
    1756 => "101101110110",
    1757 => "101101110011",
    1758 => "101101110000",
    1759 => "101101101101",
    1760 => "101101101010",
    1761 => "101101100111",
    1762 => "101101100101",
    1763 => "101101100010",
    1764 => "101101011111",
    1765 => "101101011100",
    1766 => "101101011001",
    1767 => "101101010110",
    1768 => "101101010100",
    1769 => "101101010001",
    1770 => "101101001110",
    1771 => "101101001011",
    1772 => "101101001000",
    1773 => "101101000101",
    1774 => "101101000010",
    1775 => "101100111111",
    1776 => "101100111101",
    1777 => "101100111010",
    1778 => "101100110111",
    1779 => "101100110100",
    1780 => "101100110001",
    1781 => "101100101110",
    1782 => "101100101011",
    1783 => "101100101000",
    1784 => "101100100110",
    1785 => "101100100011",
    1786 => "101100100000",
    1787 => "101100011101",
    1788 => "101100011010",
    1789 => "101100010111",
    1790 => "101100010100",
    1791 => "101100010001",
    1792 => "101100001110",
    1793 => "101100001100",
    1794 => "101100001001",
    1795 => "101100000110",
    1796 => "101100000011",
    1797 => "101100000000",
    1798 => "101011111101",
    1799 => "101011111010",
    1800 => "101011110111",
    1801 => "101011110100",
    1802 => "101011110001",
    1803 => "101011101110",
    1804 => "101011101011",
    1805 => "101011101001",
    1806 => "101011100110",
    1807 => "101011100011",
    1808 => "101011100000",
    1809 => "101011011101",
    1810 => "101011011010",
    1811 => "101011010111",
    1812 => "101011010100",
    1813 => "101011010001",
    1814 => "101011001110",
    1815 => "101011001011",
    1816 => "101011001000",
    1817 => "101011000101",
    1818 => "101011000010",
    1819 => "101010111111",
    1820 => "101010111100",
    1821 => "101010111010",
    1822 => "101010110111",
    1823 => "101010110100",
    1824 => "101010110001",
    1825 => "101010101110",
    1826 => "101010101011",
    1827 => "101010101000",
    1828 => "101010100101",
    1829 => "101010100010",
    1830 => "101010011111",
    1831 => "101010011100",
    1832 => "101010011001",
    1833 => "101010010110",
    1834 => "101010010011",
    1835 => "101010010000",
    1836 => "101010001101",
    1837 => "101010001010",
    1838 => "101010000111",
    1839 => "101010000100",
    1840 => "101010000001",
    1841 => "101001111110",
    1842 => "101001111011",
    1843 => "101001111000",
    1844 => "101001110101",
    1845 => "101001110010",
    1846 => "101001101111",
    1847 => "101001101100",
    1848 => "101001101001",
    1849 => "101001100110",
    1850 => "101001100011",
    1851 => "101001100000",
    1852 => "101001011101",
    1853 => "101001011010",
    1854 => "101001010111",
    1855 => "101001010100",
    1856 => "101001010001",
    1857 => "101001001110",
    1858 => "101001001011",
    1859 => "101001001000",
    1860 => "101001000101",
    1861 => "101001000010",
    1862 => "101000111111",
    1863 => "101000111100",
    1864 => "101000111001",
    1865 => "101000110110",
    1866 => "101000110011",
    1867 => "101000110000",
    1868 => "101000101101",
    1869 => "101000101010",
    1870 => "101000100111",
    1871 => "101000100100",
    1872 => "101000100001",
    1873 => "101000011110",
    1874 => "101000011011",
    1875 => "101000011000",
    1876 => "101000010101",
    1877 => "101000010010",
    1878 => "101000001111",
    1879 => "101000001100",
    1880 => "101000001001",
    1881 => "101000000110",
    1882 => "101000000011",
    1883 => "101000000000",
    1884 => "100111111101",
    1885 => "100111111010",
    1886 => "100111110111",
    1887 => "100111110011",
    1888 => "100111110000",
    1889 => "100111101101",
    1890 => "100111101010",
    1891 => "100111100111",
    1892 => "100111100100",
    1893 => "100111100001",
    1894 => "100111011110",
    1895 => "100111011011",
    1896 => "100111011000",
    1897 => "100111010101",
    1898 => "100111010010",
    1899 => "100111001111",
    1900 => "100111001100",
    1901 => "100111001001",
    1902 => "100111000110",
    1903 => "100111000011",
    1904 => "100111000000",
    1905 => "100110111100",
    1906 => "100110111001",
    1907 => "100110110110",
    1908 => "100110110011",
    1909 => "100110110000",
    1910 => "100110101101",
    1911 => "100110101010",
    1912 => "100110100111",
    1913 => "100110100100",
    1914 => "100110100001",
    1915 => "100110011110",
    1916 => "100110011011",
    1917 => "100110011000",
    1918 => "100110010101",
    1919 => "100110010001",
    1920 => "100110001110",
    1921 => "100110001011",
    1922 => "100110001000",
    1923 => "100110000101",
    1924 => "100110000010",
    1925 => "100101111111",
    1926 => "100101111100",
    1927 => "100101111001",
    1928 => "100101110110",
    1929 => "100101110011",
    1930 => "100101110000",
    1931 => "100101101100",
    1932 => "100101101001",
    1933 => "100101100110",
    1934 => "100101100011",
    1935 => "100101100000",
    1936 => "100101011101",
    1937 => "100101011010",
    1938 => "100101010111",
    1939 => "100101010100",
    1940 => "100101010001",
    1941 => "100101001110",
    1942 => "100101001010",
    1943 => "100101000111",
    1944 => "100101000100",
    1945 => "100101000001",
    1946 => "100100111110",
    1947 => "100100111011",
    1948 => "100100111000",
    1949 => "100100110101",
    1950 => "100100110010",
    1951 => "100100101110",
    1952 => "100100101011",
    1953 => "100100101000",
    1954 => "100100100101",
    1955 => "100100100010",
    1956 => "100100011111",
    1957 => "100100011100",
    1958 => "100100011001",
    1959 => "100100010110",
    1960 => "100100010011",
    1961 => "100100001111",
    1962 => "100100001100",
    1963 => "100100001001",
    1964 => "100100000110",
    1965 => "100100000011",
    1966 => "100100000000",
    1967 => "100011111101",
    1968 => "100011111010",
    1969 => "100011110110",
    1970 => "100011110011",
    1971 => "100011110000",
    1972 => "100011101101",
    1973 => "100011101010",
    1974 => "100011100111",
    1975 => "100011100100",
    1976 => "100011100001",
    1977 => "100011011110",
    1978 => "100011011010",
    1979 => "100011010111",
    1980 => "100011010100",
    1981 => "100011010001",
    1982 => "100011001110",
    1983 => "100011001011",
    1984 => "100011001000",
    1985 => "100011000101",
    1986 => "100011000001",
    1987 => "100010111110",
    1988 => "100010111011",
    1989 => "100010111000",
    1990 => "100010110101",
    1991 => "100010110010",
    1992 => "100010101111",
    1993 => "100010101100",
    1994 => "100010101000",
    1995 => "100010100101",
    1996 => "100010100010",
    1997 => "100010011111",
    1998 => "100010011100",
    1999 => "100010011001",
    2000 => "100010010110",
    2001 => "100010010010",
    2002 => "100010001111",
    2003 => "100010001100",
    2004 => "100010001001",
    2005 => "100010000110",
    2006 => "100010000011",
    2007 => "100010000000",
    2008 => "100001111101",
    2009 => "100001111001",
    2010 => "100001110110",
    2011 => "100001110011",
    2012 => "100001110000",
    2013 => "100001101101",
    2014 => "100001101010",
    2015 => "100001100111",
    2016 => "100001100011",
    2017 => "100001100000",
    2018 => "100001011101",
    2019 => "100001011010",
    2020 => "100001010111",
    2021 => "100001010100",
    2022 => "100001010001",
    2023 => "100001001101",
    2024 => "100001001010",
    2025 => "100001000111",
    2026 => "100001000100",
    2027 => "100001000001",
    2028 => "100000111110",
    2029 => "100000111011",
    2030 => "100000111000",
    2031 => "100000110100",
    2032 => "100000110001",
    2033 => "100000101110",
    2034 => "100000101011",
    2035 => "100000101000",
    2036 => "100000100101",
    2037 => "100000100010",
    2038 => "100000011110",
    2039 => "100000011011",
    2040 => "100000011000",
    2041 => "100000010101",
    2042 => "100000010010",
    2043 => "100000001111",
    2044 => "100000001100",
    2045 => "100000001000",
    2046 => "100000000101",
    2047 => "100000000010",
    2048 => "011111111111",
    2049 => "011111111100",
    2050 => "011111111001",
    2051 => "011111110110",
    2052 => "011111110010",
    2053 => "011111101111",
    2054 => "011111101100",
    2055 => "011111101001",
    2056 => "011111100110",
    2057 => "011111100011",
    2058 => "011111100000",
    2059 => "011111011100",
    2060 => "011111011001",
    2061 => "011111010110",
    2062 => "011111010011",
    2063 => "011111010000",
    2064 => "011111001101",
    2065 => "011111001010",
    2066 => "011111000110",
    2067 => "011111000011",
    2068 => "011111000000",
    2069 => "011110111101",
    2070 => "011110111010",
    2071 => "011110110111",
    2072 => "011110110100",
    2073 => "011110110001",
    2074 => "011110101101",
    2075 => "011110101010",
    2076 => "011110100111",
    2077 => "011110100100",
    2078 => "011110100001",
    2079 => "011110011110",
    2080 => "011110011011",
    2081 => "011110010111",
    2082 => "011110010100",
    2083 => "011110010001",
    2084 => "011110001110",
    2085 => "011110001011",
    2086 => "011110001000",
    2087 => "011110000101",
    2088 => "011110000001",
    2089 => "011101111110",
    2090 => "011101111011",
    2091 => "011101111000",
    2092 => "011101110101",
    2093 => "011101110010",
    2094 => "011101101111",
    2095 => "011101101100",
    2096 => "011101101000",
    2097 => "011101100101",
    2098 => "011101100010",
    2099 => "011101011111",
    2100 => "011101011100",
    2101 => "011101011001",
    2102 => "011101010110",
    2103 => "011101010010",
    2104 => "011101001111",
    2105 => "011101001100",
    2106 => "011101001001",
    2107 => "011101000110",
    2108 => "011101000011",
    2109 => "011101000000",
    2110 => "011100111101",
    2111 => "011100111001",
    2112 => "011100110110",
    2113 => "011100110011",
    2114 => "011100110000",
    2115 => "011100101101",
    2116 => "011100101010",
    2117 => "011100100111",
    2118 => "011100100100",
    2119 => "011100100000",
    2120 => "011100011101",
    2121 => "011100011010",
    2122 => "011100010111",
    2123 => "011100010100",
    2124 => "011100010001",
    2125 => "011100001110",
    2126 => "011100001011",
    2127 => "011100001000",
    2128 => "011100000100",
    2129 => "011100000001",
    2130 => "011011111110",
    2131 => "011011111011",
    2132 => "011011111000",
    2133 => "011011110101",
    2134 => "011011110010",
    2135 => "011011101111",
    2136 => "011011101011",
    2137 => "011011101000",
    2138 => "011011100101",
    2139 => "011011100010",
    2140 => "011011011111",
    2141 => "011011011100",
    2142 => "011011011001",
    2143 => "011011010110",
    2144 => "011011010011",
    2145 => "011011010000",
    2146 => "011011001100",
    2147 => "011011001001",
    2148 => "011011000110",
    2149 => "011011000011",
    2150 => "011011000000",
    2151 => "011010111101",
    2152 => "011010111010",
    2153 => "011010110111",
    2154 => "011010110100",
    2155 => "011010110000",
    2156 => "011010101101",
    2157 => "011010101010",
    2158 => "011010100111",
    2159 => "011010100100",
    2160 => "011010100001",
    2161 => "011010011110",
    2162 => "011010011011",
    2163 => "011010011000",
    2164 => "011010010101",
    2165 => "011010010010",
    2166 => "011010001110",
    2167 => "011010001011",
    2168 => "011010001000",
    2169 => "011010000101",
    2170 => "011010000010",
    2171 => "011001111111",
    2172 => "011001111100",
    2173 => "011001111001",
    2174 => "011001110110",
    2175 => "011001110011",
    2176 => "011001110000",
    2177 => "011001101101",
    2178 => "011001101001",
    2179 => "011001100110",
    2180 => "011001100011",
    2181 => "011001100000",
    2182 => "011001011101",
    2183 => "011001011010",
    2184 => "011001010111",
    2185 => "011001010100",
    2186 => "011001010001",
    2187 => "011001001110",
    2188 => "011001001011",
    2189 => "011001001000",
    2190 => "011001000101",
    2191 => "011001000010",
    2192 => "011000111110",
    2193 => "011000111011",
    2194 => "011000111000",
    2195 => "011000110101",
    2196 => "011000110010",
    2197 => "011000101111",
    2198 => "011000101100",
    2199 => "011000101001",
    2200 => "011000100110",
    2201 => "011000100011",
    2202 => "011000100000",
    2203 => "011000011101",
    2204 => "011000011010",
    2205 => "011000010111",
    2206 => "011000010100",
    2207 => "011000010001",
    2208 => "011000001110",
    2209 => "011000001011",
    2210 => "011000000111",
    2211 => "011000000100",
    2212 => "011000000001",
    2213 => "010111111110",
    2214 => "010111111011",
    2215 => "010111111000",
    2216 => "010111110101",
    2217 => "010111110010",
    2218 => "010111101111",
    2219 => "010111101100",
    2220 => "010111101001",
    2221 => "010111100110",
    2222 => "010111100011",
    2223 => "010111100000",
    2224 => "010111011101",
    2225 => "010111011010",
    2226 => "010111010111",
    2227 => "010111010100",
    2228 => "010111010001",
    2229 => "010111001110",
    2230 => "010111001011",
    2231 => "010111001000",
    2232 => "010111000101",
    2233 => "010111000010",
    2234 => "010110111111",
    2235 => "010110111100",
    2236 => "010110111001",
    2237 => "010110110110",
    2238 => "010110110011",
    2239 => "010110110000",
    2240 => "010110101101",
    2241 => "010110101010",
    2242 => "010110100111",
    2243 => "010110100100",
    2244 => "010110100001",
    2245 => "010110011110",
    2246 => "010110011011",
    2247 => "010110011000",
    2248 => "010110010101",
    2249 => "010110010010",
    2250 => "010110001111",
    2251 => "010110001100",
    2252 => "010110001001",
    2253 => "010110000110",
    2254 => "010110000011",
    2255 => "010110000000",
    2256 => "010101111101",
    2257 => "010101111010",
    2258 => "010101110111",
    2259 => "010101110100",
    2260 => "010101110001",
    2261 => "010101101110",
    2262 => "010101101011",
    2263 => "010101101000",
    2264 => "010101100101",
    2265 => "010101100010",
    2266 => "010101011111",
    2267 => "010101011100",
    2268 => "010101011001",
    2269 => "010101010110",
    2270 => "010101010011",
    2271 => "010101010000",
    2272 => "010101001101",
    2273 => "010101001010",
    2274 => "010101000111",
    2275 => "010101000100",
    2276 => "010101000010",
    2277 => "010100111111",
    2278 => "010100111100",
    2279 => "010100111001",
    2280 => "010100110110",
    2281 => "010100110011",
    2282 => "010100110000",
    2283 => "010100101101",
    2284 => "010100101010",
    2285 => "010100100111",
    2286 => "010100100100",
    2287 => "010100100001",
    2288 => "010100011110",
    2289 => "010100011011",
    2290 => "010100011000",
    2291 => "010100010101",
    2292 => "010100010011",
    2293 => "010100010000",
    2294 => "010100001101",
    2295 => "010100001010",
    2296 => "010100000111",
    2297 => "010100000100",
    2298 => "010100000001",
    2299 => "010011111110",
    2300 => "010011111011",
    2301 => "010011111000",
    2302 => "010011110101",
    2303 => "010011110010",
    2304 => "010011110000",
    2305 => "010011101101",
    2306 => "010011101010",
    2307 => "010011100111",
    2308 => "010011100100",
    2309 => "010011100001",
    2310 => "010011011110",
    2311 => "010011011011",
    2312 => "010011011000",
    2313 => "010011010110",
    2314 => "010011010011",
    2315 => "010011010000",
    2316 => "010011001101",
    2317 => "010011001010",
    2318 => "010011000111",
    2319 => "010011000100",
    2320 => "010011000001",
    2321 => "010010111111",
    2322 => "010010111100",
    2323 => "010010111001",
    2324 => "010010110110",
    2325 => "010010110011",
    2326 => "010010110000",
    2327 => "010010101101",
    2328 => "010010101010",
    2329 => "010010101000",
    2330 => "010010100101",
    2331 => "010010100010",
    2332 => "010010011111",
    2333 => "010010011100",
    2334 => "010010011001",
    2335 => "010010010111",
    2336 => "010010010100",
    2337 => "010010010001",
    2338 => "010010001110",
    2339 => "010010001011",
    2340 => "010010001000",
    2341 => "010010000110",
    2342 => "010010000011",
    2343 => "010010000000",
    2344 => "010001111101",
    2345 => "010001111010",
    2346 => "010001110111",
    2347 => "010001110101",
    2348 => "010001110010",
    2349 => "010001101111",
    2350 => "010001101100",
    2351 => "010001101001",
    2352 => "010001100111",
    2353 => "010001100100",
    2354 => "010001100001",
    2355 => "010001011110",
    2356 => "010001011011",
    2357 => "010001011001",
    2358 => "010001010110",
    2359 => "010001010011",
    2360 => "010001010000",
    2361 => "010001001101",
    2362 => "010001001011",
    2363 => "010001001000",
    2364 => "010001000101",
    2365 => "010001000010",
    2366 => "010001000000",
    2367 => "010000111101",
    2368 => "010000111010",
    2369 => "010000110111",
    2370 => "010000110100",
    2371 => "010000110010",
    2372 => "010000101111",
    2373 => "010000101100",
    2374 => "010000101001",
    2375 => "010000100111",
    2376 => "010000100100",
    2377 => "010000100001",
    2378 => "010000011110",
    2379 => "010000011100",
    2380 => "010000011001",
    2381 => "010000010110",
    2382 => "010000010011",
    2383 => "010000010001",
    2384 => "010000001110",
    2385 => "010000001011",
    2386 => "010000001000",
    2387 => "010000000110",
    2388 => "010000000011",
    2389 => "010000000000",
    2390 => "001111111110",
    2391 => "001111111011",
    2392 => "001111111000",
    2393 => "001111110101",
    2394 => "001111110011",
    2395 => "001111110000",
    2396 => "001111101101",
    2397 => "001111101011",
    2398 => "001111101000",
    2399 => "001111100101",
    2400 => "001111100011",
    2401 => "001111100000",
    2402 => "001111011101",
    2403 => "001111011010",
    2404 => "001111011000",
    2405 => "001111010101",
    2406 => "001111010010",
    2407 => "001111010000",
    2408 => "001111001101",
    2409 => "001111001010",
    2410 => "001111001000",
    2411 => "001111000101",
    2412 => "001111000010",
    2413 => "001111000000",
    2414 => "001110111101",
    2415 => "001110111010",
    2416 => "001110111000",
    2417 => "001110110101",
    2418 => "001110110010",
    2419 => "001110110000",
    2420 => "001110101101",
    2421 => "001110101011",
    2422 => "001110101000",
    2423 => "001110100101",
    2424 => "001110100011",
    2425 => "001110100000",
    2426 => "001110011101",
    2427 => "001110011011",
    2428 => "001110011000",
    2429 => "001110010101",
    2430 => "001110010011",
    2431 => "001110010000",
    2432 => "001110001110",
    2433 => "001110001011",
    2434 => "001110001000",
    2435 => "001110000110",
    2436 => "001110000011",
    2437 => "001110000001",
    2438 => "001101111110",
    2439 => "001101111011",
    2440 => "001101111001",
    2441 => "001101110110",
    2442 => "001101110100",
    2443 => "001101110001",
    2444 => "001101101111",
    2445 => "001101101100",
    2446 => "001101101001",
    2447 => "001101100111",
    2448 => "001101100100",
    2449 => "001101100010",
    2450 => "001101011111",
    2451 => "001101011101",
    2452 => "001101011010",
    2453 => "001101010111",
    2454 => "001101010101",
    2455 => "001101010010",
    2456 => "001101010000",
    2457 => "001101001101",
    2458 => "001101001011",
    2459 => "001101001000",
    2460 => "001101000110",
    2461 => "001101000011",
    2462 => "001101000001",
    2463 => "001100111110",
    2464 => "001100111011",
    2465 => "001100111001",
    2466 => "001100110110",
    2467 => "001100110100",
    2468 => "001100110001",
    2469 => "001100101111",
    2470 => "001100101100",
    2471 => "001100101010",
    2472 => "001100100111",
    2473 => "001100100101",
    2474 => "001100100010",
    2475 => "001100100000",
    2476 => "001100011101",
    2477 => "001100011011",
    2478 => "001100011000",
    2479 => "001100010110",
    2480 => "001100010100",
    2481 => "001100010001",
    2482 => "001100001111",
    2483 => "001100001100",
    2484 => "001100001010",
    2485 => "001100000111",
    2486 => "001100000101",
    2487 => "001100000010",
    2488 => "001100000000",
    2489 => "001011111101",
    2490 => "001011111011",
    2491 => "001011111000",
    2492 => "001011110110",
    2493 => "001011110100",
    2494 => "001011110001",
    2495 => "001011101111",
    2496 => "001011101100",
    2497 => "001011101010",
    2498 => "001011100111",
    2499 => "001011100101",
    2500 => "001011100011",
    2501 => "001011100000",
    2502 => "001011011110",
    2503 => "001011011011",
    2504 => "001011011001",
    2505 => "001011010111",
    2506 => "001011010100",
    2507 => "001011010010",
    2508 => "001011001111",
    2509 => "001011001101",
    2510 => "001011001011",
    2511 => "001011001000",
    2512 => "001011000110",
    2513 => "001011000011",
    2514 => "001011000001",
    2515 => "001010111111",
    2516 => "001010111100",
    2517 => "001010111010",
    2518 => "001010111000",
    2519 => "001010110101",
    2520 => "001010110011",
    2521 => "001010110001",
    2522 => "001010101110",
    2523 => "001010101100",
    2524 => "001010101010",
    2525 => "001010100111",
    2526 => "001010100101",
    2527 => "001010100011",
    2528 => "001010100000",
    2529 => "001010011110",
    2530 => "001010011100",
    2531 => "001010011001",
    2532 => "001010010111",
    2533 => "001010010101",
    2534 => "001010010010",
    2535 => "001010010000",
    2536 => "001010001110",
    2537 => "001010001011",
    2538 => "001010001001",
    2539 => "001010000111",
    2540 => "001010000101",
    2541 => "001010000010",
    2542 => "001010000000",
    2543 => "001001111110",
    2544 => "001001111011",
    2545 => "001001111001",
    2546 => "001001110111",
    2547 => "001001110101",
    2548 => "001001110010",
    2549 => "001001110000",
    2550 => "001001101110",
    2551 => "001001101100",
    2552 => "001001101001",
    2553 => "001001100111",
    2554 => "001001100101",
    2555 => "001001100011",
    2556 => "001001100000",
    2557 => "001001011110",
    2558 => "001001011100",
    2559 => "001001011010",
    2560 => "001001010111",
    2561 => "001001010101",
    2562 => "001001010011",
    2563 => "001001010001",
    2564 => "001001001111",
    2565 => "001001001100",
    2566 => "001001001010",
    2567 => "001001001000",
    2568 => "001001000110",
    2569 => "001001000100",
    2570 => "001001000001",
    2571 => "001000111111",
    2572 => "001000111101",
    2573 => "001000111011",
    2574 => "001000111001",
    2575 => "001000110111",
    2576 => "001000110100",
    2577 => "001000110010",
    2578 => "001000110000",
    2579 => "001000101110",
    2580 => "001000101100",
    2581 => "001000101010",
    2582 => "001000100111",
    2583 => "001000100101",
    2584 => "001000100011",
    2585 => "001000100001",
    2586 => "001000011111",
    2587 => "001000011101",
    2588 => "001000011011",
    2589 => "001000011000",
    2590 => "001000010110",
    2591 => "001000010100",
    2592 => "001000010010",
    2593 => "001000010000",
    2594 => "001000001110",
    2595 => "001000001100",
    2596 => "001000001010",
    2597 => "001000001000",
    2598 => "001000000110",
    2599 => "001000000011",
    2600 => "001000000001",
    2601 => "000111111111",
    2602 => "000111111101",
    2603 => "000111111011",
    2604 => "000111111001",
    2605 => "000111110111",
    2606 => "000111110101",
    2607 => "000111110011",
    2608 => "000111110001",
    2609 => "000111101111",
    2610 => "000111101101",
    2611 => "000111101011",
    2612 => "000111101001",
    2613 => "000111100111",
    2614 => "000111100101",
    2615 => "000111100011",
    2616 => "000111100001",
    2617 => "000111011111",
    2618 => "000111011101",
    2619 => "000111011011",
    2620 => "000111011001",
    2621 => "000111010111",
    2622 => "000111010100",
    2623 => "000111010011",
    2624 => "000111010001",
    2625 => "000111001111",
    2626 => "000111001101",
    2627 => "000111001011",
    2628 => "000111001001",
    2629 => "000111000111",
    2630 => "000111000101",
    2631 => "000111000011",
    2632 => "000111000001",
    2633 => "000110111111",
    2634 => "000110111101",
    2635 => "000110111011",
    2636 => "000110111001",
    2637 => "000110110111",
    2638 => "000110110101",
    2639 => "000110110011",
    2640 => "000110110001",
    2641 => "000110101111",
    2642 => "000110101101",
    2643 => "000110101011",
    2644 => "000110101001",
    2645 => "000110100111",
    2646 => "000110100110",
    2647 => "000110100100",
    2648 => "000110100010",
    2649 => "000110100000",
    2650 => "000110011110",
    2651 => "000110011100",
    2652 => "000110011010",
    2653 => "000110011000",
    2654 => "000110010110",
    2655 => "000110010101",
    2656 => "000110010011",
    2657 => "000110010001",
    2658 => "000110001111",
    2659 => "000110001101",
    2660 => "000110001011",
    2661 => "000110001001",
    2662 => "000110001000",
    2663 => "000110000110",
    2664 => "000110000100",
    2665 => "000110000010",
    2666 => "000110000000",
    2667 => "000101111110",
    2668 => "000101111101",
    2669 => "000101111011",
    2670 => "000101111001",
    2671 => "000101110111",
    2672 => "000101110101",
    2673 => "000101110011",
    2674 => "000101110010",
    2675 => "000101110000",
    2676 => "000101101110",
    2677 => "000101101100",
    2678 => "000101101010",
    2679 => "000101101001",
    2680 => "000101100111",
    2681 => "000101100101",
    2682 => "000101100011",
    2683 => "000101100010",
    2684 => "000101100000",
    2685 => "000101011110",
    2686 => "000101011100",
    2687 => "000101011011",
    2688 => "000101011001",
    2689 => "000101010111",
    2690 => "000101010101",
    2691 => "000101010100",
    2692 => "000101010010",
    2693 => "000101010000",
    2694 => "000101001110",
    2695 => "000101001101",
    2696 => "000101001011",
    2697 => "000101001001",
    2698 => "000101001000",
    2699 => "000101000110",
    2700 => "000101000100",
    2701 => "000101000010",
    2702 => "000101000001",
    2703 => "000100111111",
    2704 => "000100111101",
    2705 => "000100111100",
    2706 => "000100111010",
    2707 => "000100111000",
    2708 => "000100110111",
    2709 => "000100110101",
    2710 => "000100110011",
    2711 => "000100110010",
    2712 => "000100110000",
    2713 => "000100101110",
    2714 => "000100101101",
    2715 => "000100101011",
    2716 => "000100101010",
    2717 => "000100101000",
    2718 => "000100100110",
    2719 => "000100100101",
    2720 => "000100100011",
    2721 => "000100100001",
    2722 => "000100100000",
    2723 => "000100011110",
    2724 => "000100011101",
    2725 => "000100011011",
    2726 => "000100011001",
    2727 => "000100011000",
    2728 => "000100010110",
    2729 => "000100010101",
    2730 => "000100010011",
    2731 => "000100010010",
    2732 => "000100010000",
    2733 => "000100001110",
    2734 => "000100001101",
    2735 => "000100001011",
    2736 => "000100001010",
    2737 => "000100001000",
    2738 => "000100000111",
    2739 => "000100000101",
    2740 => "000100000100",
    2741 => "000100000010",
    2742 => "000100000001",
    2743 => "000011111111",
    2744 => "000011111110",
    2745 => "000011111100",
    2746 => "000011111011",
    2747 => "000011111001",
    2748 => "000011111000",
    2749 => "000011110110",
    2750 => "000011110101",
    2751 => "000011110011",
    2752 => "000011110010",
    2753 => "000011110000",
    2754 => "000011101111",
    2755 => "000011101101",
    2756 => "000011101100",
    2757 => "000011101010",
    2758 => "000011101001",
    2759 => "000011100111",
    2760 => "000011100110",
    2761 => "000011100100",
    2762 => "000011100011",
    2763 => "000011100010",
    2764 => "000011100000",
    2765 => "000011011111",
    2766 => "000011011101",
    2767 => "000011011100",
    2768 => "000011011010",
    2769 => "000011011001",
    2770 => "000011011000",
    2771 => "000011010110",
    2772 => "000011010101",
    2773 => "000011010011",
    2774 => "000011010010",
    2775 => "000011010001",
    2776 => "000011001111",
    2777 => "000011001110",
    2778 => "000011001101",
    2779 => "000011001011",
    2780 => "000011001010",
    2781 => "000011001000",
    2782 => "000011000111",
    2783 => "000011000110",
    2784 => "000011000100",
    2785 => "000011000011",
    2786 => "000011000010",
    2787 => "000011000000",
    2788 => "000010111111",
    2789 => "000010111110",
    2790 => "000010111100",
    2791 => "000010111011",
    2792 => "000010111010",
    2793 => "000010111000",
    2794 => "000010110111",
    2795 => "000010110110",
    2796 => "000010110101",
    2797 => "000010110011",
    2798 => "000010110010",
    2799 => "000010110001",
    2800 => "000010101111",
    2801 => "000010101110",
    2802 => "000010101101",
    2803 => "000010101100",
    2804 => "000010101010",
    2805 => "000010101001",
    2806 => "000010101000",
    2807 => "000010100111",
    2808 => "000010100101",
    2809 => "000010100100",
    2810 => "000010100011",
    2811 => "000010100010",
    2812 => "000010100000",
    2813 => "000010011111",
    2814 => "000010011110",
    2815 => "000010011101",
    2816 => "000010011100",
    2817 => "000010011010",
    2818 => "000010011001",
    2819 => "000010011000",
    2820 => "000010010111",
    2821 => "000010010110",
    2822 => "000010010101",
    2823 => "000010010011",
    2824 => "000010010010",
    2825 => "000010010001",
    2826 => "000010010000",
    2827 => "000010001111",
    2828 => "000010001110",
    2829 => "000010001100",
    2830 => "000010001011",
    2831 => "000010001010",
    2832 => "000010001001",
    2833 => "000010001000",
    2834 => "000010000111",
    2835 => "000010000110",
    2836 => "000010000101",
    2837 => "000010000011",
    2838 => "000010000010",
    2839 => "000010000001",
    2840 => "000010000000",
    2841 => "000001111111",
    2842 => "000001111110",
    2843 => "000001111101",
    2844 => "000001111100",
    2845 => "000001111011",
    2846 => "000001111010",
    2847 => "000001111001",
    2848 => "000001110111",
    2849 => "000001110110",
    2850 => "000001110101",
    2851 => "000001110100",
    2852 => "000001110011",
    2853 => "000001110010",
    2854 => "000001110001",
    2855 => "000001110000",
    2856 => "000001101111",
    2857 => "000001101110",
    2858 => "000001101101",
    2859 => "000001101100",
    2860 => "000001101011",
    2861 => "000001101010",
    2862 => "000001101001",
    2863 => "000001101000",
    2864 => "000001100111",
    2865 => "000001100110",
    2866 => "000001100101",
    2867 => "000001100100",
    2868 => "000001100011",
    2869 => "000001100010",
    2870 => "000001100001",
    2871 => "000001100000",
    2872 => "000001011111",
    2873 => "000001011110",
    2874 => "000001011110",
    2875 => "000001011101",
    2876 => "000001011100",
    2877 => "000001011011",
    2878 => "000001011010",
    2879 => "000001011001",
    2880 => "000001011000",
    2881 => "000001010111",
    2882 => "000001010110",
    2883 => "000001010101",
    2884 => "000001010100",
    2885 => "000001010011",
    2886 => "000001010011",
    2887 => "000001010010",
    2888 => "000001010001",
    2889 => "000001010000",
    2890 => "000001001111",
    2891 => "000001001110",
    2892 => "000001001101",
    2893 => "000001001101",
    2894 => "000001001100",
    2895 => "000001001011",
    2896 => "000001001010",
    2897 => "000001001001",
    2898 => "000001001000",
    2899 => "000001000111",
    2900 => "000001000111",
    2901 => "000001000110",
    2902 => "000001000101",
    2903 => "000001000100",
    2904 => "000001000011",
    2905 => "000001000011",
    2906 => "000001000010",
    2907 => "000001000001",
    2908 => "000001000000",
    2909 => "000000111111",
    2910 => "000000111111",
    2911 => "000000111110",
    2912 => "000000111101",
    2913 => "000000111100",
    2914 => "000000111100",
    2915 => "000000111011",
    2916 => "000000111010",
    2917 => "000000111001",
    2918 => "000000111001",
    2919 => "000000111000",
    2920 => "000000110111",
    2921 => "000000110110",
    2922 => "000000110110",
    2923 => "000000110101",
    2924 => "000000110100",
    2925 => "000000110100",
    2926 => "000000110011",
    2927 => "000000110010",
    2928 => "000000110010",
    2929 => "000000110001",
    2930 => "000000110000",
    2931 => "000000110000",
    2932 => "000000101111",
    2933 => "000000101110",
    2934 => "000000101110",
    2935 => "000000101101",
    2936 => "000000101100",
    2937 => "000000101100",
    2938 => "000000101011",
    2939 => "000000101010",
    2940 => "000000101010",
    2941 => "000000101001",
    2942 => "000000101000",
    2943 => "000000101000",
    2944 => "000000100111",
    2945 => "000000100111",
    2946 => "000000100110",
    2947 => "000000100101",
    2948 => "000000100101",
    2949 => "000000100100",
    2950 => "000000100100",
    2951 => "000000100011",
    2952 => "000000100010",
    2953 => "000000100010",
    2954 => "000000100001",
    2955 => "000000100001",
    2956 => "000000100000",
    2957 => "000000100000",
    2958 => "000000011111",
    2959 => "000000011110",
    2960 => "000000011110",
    2961 => "000000011101",
    2962 => "000000011101",
    2963 => "000000011100",
    2964 => "000000011100",
    2965 => "000000011011",
    2966 => "000000011011",
    2967 => "000000011010",
    2968 => "000000011010",
    2969 => "000000011001",
    2970 => "000000011001",
    2971 => "000000011000",
    2972 => "000000011000",
    2973 => "000000010111",
    2974 => "000000010111",
    2975 => "000000010110",
    2976 => "000000010110",
    2977 => "000000010110",
    2978 => "000000010101",
    2979 => "000000010101",
    2980 => "000000010100",
    2981 => "000000010100",
    2982 => "000000010011",
    2983 => "000000010011",
    2984 => "000000010010",
    2985 => "000000010010",
    2986 => "000000010010",
    2987 => "000000010001",
    2988 => "000000010001",
    2989 => "000000010000",
    2990 => "000000010000",
    2991 => "000000010000",
    2992 => "000000001111",
    2993 => "000000001111",
    2994 => "000000001110",
    2995 => "000000001110",
    2996 => "000000001110",
    2997 => "000000001101",
    2998 => "000000001101",
    2999 => "000000001101",
    3000 => "000000001100",
    3001 => "000000001100",
    3002 => "000000001100",
    3003 => "000000001011",
    3004 => "000000001011",
    3005 => "000000001011",
    3006 => "000000001010",
    3007 => "000000001010",
    3008 => "000000001010",
    3009 => "000000001001",
    3010 => "000000001001",
    3011 => "000000001001",
    3012 => "000000001000",
    3013 => "000000001000",
    3014 => "000000001000",
    3015 => "000000001000",
    3016 => "000000000111",
    3017 => "000000000111",
    3018 => "000000000111",
    3019 => "000000000111",
    3020 => "000000000110",
    3021 => "000000000110",
    3022 => "000000000110",
    3023 => "000000000110",
    3024 => "000000000101",
    3025 => "000000000101",
    3026 => "000000000101",
    3027 => "000000000101",
    3028 => "000000000100",
    3029 => "000000000100",
    3030 => "000000000100",
    3031 => "000000000100",
    3032 => "000000000100",
    3033 => "000000000011",
    3034 => "000000000011",
    3035 => "000000000011",
    3036 => "000000000011",
    3037 => "000000000011",
    3038 => "000000000011",
    3039 => "000000000010",
    3040 => "000000000010",
    3041 => "000000000010",
    3042 => "000000000010",
    3043 => "000000000010",
    3044 => "000000000010",
    3045 => "000000000010",
    3046 => "000000000001",
    3047 => "000000000001",
    3048 => "000000000001",
    3049 => "000000000001",
    3050 => "000000000001",
    3051 => "000000000001",
    3052 => "000000000001",
    3053 => "000000000001",
    3054 => "000000000001",
    3055 => "000000000001",
    3056 => "000000000000",
    3057 => "000000000000",
    3058 => "000000000000",
    3059 => "000000000000",
    3060 => "000000000000",
    3061 => "000000000000",
    3062 => "000000000000",
    3063 => "000000000000",
    3064 => "000000000000",
    3065 => "000000000000",
    3066 => "000000000000",
    3067 => "000000000000",
    3068 => "000000000000",
    3069 => "000000000000",
    3070 => "000000000000",
    3071 => "000000000000",
    3072 => "000000000000",
    3073 => "000000000000",
    3074 => "000000000000",
    3075 => "000000000000",
    3076 => "000000000000",
    3077 => "000000000000",
    3078 => "000000000000",
    3079 => "000000000000",
    3080 => "000000000000",
    3081 => "000000000000",
    3082 => "000000000000",
    3083 => "000000000000",
    3084 => "000000000000",
    3085 => "000000000000",
    3086 => "000000000000",
    3087 => "000000000000",
    3088 => "000000000000",
    3089 => "000000000001",
    3090 => "000000000001",
    3091 => "000000000001",
    3092 => "000000000001",
    3093 => "000000000001",
    3094 => "000000000001",
    3095 => "000000000001",
    3096 => "000000000001",
    3097 => "000000000001",
    3098 => "000000000001",
    3099 => "000000000010",
    3100 => "000000000010",
    3101 => "000000000010",
    3102 => "000000000010",
    3103 => "000000000010",
    3104 => "000000000010",
    3105 => "000000000010",
    3106 => "000000000011",
    3107 => "000000000011",
    3108 => "000000000011",
    3109 => "000000000011",
    3110 => "000000000011",
    3111 => "000000000011",
    3112 => "000000000100",
    3113 => "000000000100",
    3114 => "000000000100",
    3115 => "000000000100",
    3116 => "000000000100",
    3117 => "000000000101",
    3118 => "000000000101",
    3119 => "000000000101",
    3120 => "000000000101",
    3121 => "000000000110",
    3122 => "000000000110",
    3123 => "000000000110",
    3124 => "000000000110",
    3125 => "000000000111",
    3126 => "000000000111",
    3127 => "000000000111",
    3128 => "000000000111",
    3129 => "000000001000",
    3130 => "000000001000",
    3131 => "000000001000",
    3132 => "000000001000",
    3133 => "000000001001",
    3134 => "000000001001",
    3135 => "000000001001",
    3136 => "000000001010",
    3137 => "000000001010",
    3138 => "000000001010",
    3139 => "000000001011",
    3140 => "000000001011",
    3141 => "000000001011",
    3142 => "000000001100",
    3143 => "000000001100",
    3144 => "000000001100",
    3145 => "000000001101",
    3146 => "000000001101",
    3147 => "000000001101",
    3148 => "000000001110",
    3149 => "000000001110",
    3150 => "000000001110",
    3151 => "000000001111",
    3152 => "000000001111",
    3153 => "000000010000",
    3154 => "000000010000",
    3155 => "000000010000",
    3156 => "000000010001",
    3157 => "000000010001",
    3158 => "000000010010",
    3159 => "000000010010",
    3160 => "000000010010",
    3161 => "000000010011",
    3162 => "000000010011",
    3163 => "000000010100",
    3164 => "000000010100",
    3165 => "000000010101",
    3166 => "000000010101",
    3167 => "000000010110",
    3168 => "000000010110",
    3169 => "000000010110",
    3170 => "000000010111",
    3171 => "000000010111",
    3172 => "000000011000",
    3173 => "000000011000",
    3174 => "000000011001",
    3175 => "000000011001",
    3176 => "000000011010",
    3177 => "000000011010",
    3178 => "000000011011",
    3179 => "000000011011",
    3180 => "000000011100",
    3181 => "000000011100",
    3182 => "000000011101",
    3183 => "000000011101",
    3184 => "000000011110",
    3185 => "000000011110",
    3186 => "000000011111",
    3187 => "000000100000",
    3188 => "000000100000",
    3189 => "000000100001",
    3190 => "000000100001",
    3191 => "000000100010",
    3192 => "000000100010",
    3193 => "000000100011",
    3194 => "000000100100",
    3195 => "000000100100",
    3196 => "000000100101",
    3197 => "000000100101",
    3198 => "000000100110",
    3199 => "000000100111",
    3200 => "000000100111",
    3201 => "000000101000",
    3202 => "000000101000",
    3203 => "000000101001",
    3204 => "000000101010",
    3205 => "000000101010",
    3206 => "000000101011",
    3207 => "000000101100",
    3208 => "000000101100",
    3209 => "000000101101",
    3210 => "000000101110",
    3211 => "000000101110",
    3212 => "000000101111",
    3213 => "000000110000",
    3214 => "000000110000",
    3215 => "000000110001",
    3216 => "000000110010",
    3217 => "000000110010",
    3218 => "000000110011",
    3219 => "000000110100",
    3220 => "000000110100",
    3221 => "000000110101",
    3222 => "000000110110",
    3223 => "000000110110",
    3224 => "000000110111",
    3225 => "000000111000",
    3226 => "000000111001",
    3227 => "000000111001",
    3228 => "000000111010",
    3229 => "000000111011",
    3230 => "000000111100",
    3231 => "000000111100",
    3232 => "000000111101",
    3233 => "000000111110",
    3234 => "000000111111",
    3235 => "000000111111",
    3236 => "000001000000",
    3237 => "000001000001",
    3238 => "000001000010",
    3239 => "000001000011",
    3240 => "000001000011",
    3241 => "000001000100",
    3242 => "000001000101",
    3243 => "000001000110",
    3244 => "000001000111",
    3245 => "000001000111",
    3246 => "000001001000",
    3247 => "000001001001",
    3248 => "000001001010",
    3249 => "000001001011",
    3250 => "000001001100",
    3251 => "000001001101",
    3252 => "000001001101",
    3253 => "000001001110",
    3254 => "000001001111",
    3255 => "000001010000",
    3256 => "000001010001",
    3257 => "000001010010",
    3258 => "000001010011",
    3259 => "000001010011",
    3260 => "000001010100",
    3261 => "000001010101",
    3262 => "000001010110",
    3263 => "000001010111",
    3264 => "000001011000",
    3265 => "000001011001",
    3266 => "000001011010",
    3267 => "000001011011",
    3268 => "000001011100",
    3269 => "000001011101",
    3270 => "000001011110",
    3271 => "000001011110",
    3272 => "000001011111",
    3273 => "000001100000",
    3274 => "000001100001",
    3275 => "000001100010",
    3276 => "000001100011",
    3277 => "000001100100",
    3278 => "000001100101",
    3279 => "000001100110",
    3280 => "000001100111",
    3281 => "000001101000",
    3282 => "000001101001",
    3283 => "000001101010",
    3284 => "000001101011",
    3285 => "000001101100",
    3286 => "000001101101",
    3287 => "000001101110",
    3288 => "000001101111",
    3289 => "000001110000",
    3290 => "000001110001",
    3291 => "000001110010",
    3292 => "000001110011",
    3293 => "000001110100",
    3294 => "000001110101",
    3295 => "000001110110",
    3296 => "000001110111",
    3297 => "000001111001",
    3298 => "000001111010",
    3299 => "000001111011",
    3300 => "000001111100",
    3301 => "000001111101",
    3302 => "000001111110",
    3303 => "000001111111",
    3304 => "000010000000",
    3305 => "000010000001",
    3306 => "000010000010",
    3307 => "000010000011",
    3308 => "000010000101",
    3309 => "000010000110",
    3310 => "000010000111",
    3311 => "000010001000",
    3312 => "000010001001",
    3313 => "000010001010",
    3314 => "000010001011",
    3315 => "000010001100",
    3316 => "000010001110",
    3317 => "000010001111",
    3318 => "000010010000",
    3319 => "000010010001",
    3320 => "000010010010",
    3321 => "000010010011",
    3322 => "000010010101",
    3323 => "000010010110",
    3324 => "000010010111",
    3325 => "000010011000",
    3326 => "000010011001",
    3327 => "000010011010",
    3328 => "000010011100",
    3329 => "000010011101",
    3330 => "000010011110",
    3331 => "000010011111",
    3332 => "000010100000",
    3333 => "000010100010",
    3334 => "000010100011",
    3335 => "000010100100",
    3336 => "000010100101",
    3337 => "000010100111",
    3338 => "000010101000",
    3339 => "000010101001",
    3340 => "000010101010",
    3341 => "000010101100",
    3342 => "000010101101",
    3343 => "000010101110",
    3344 => "000010101111",
    3345 => "000010110001",
    3346 => "000010110010",
    3347 => "000010110011",
    3348 => "000010110101",
    3349 => "000010110110",
    3350 => "000010110111",
    3351 => "000010111000",
    3352 => "000010111010",
    3353 => "000010111011",
    3354 => "000010111100",
    3355 => "000010111110",
    3356 => "000010111111",
    3357 => "000011000000",
    3358 => "000011000010",
    3359 => "000011000011",
    3360 => "000011000100",
    3361 => "000011000110",
    3362 => "000011000111",
    3363 => "000011001000",
    3364 => "000011001010",
    3365 => "000011001011",
    3366 => "000011001101",
    3367 => "000011001110",
    3368 => "000011001111",
    3369 => "000011010001",
    3370 => "000011010010",
    3371 => "000011010011",
    3372 => "000011010101",
    3373 => "000011010110",
    3374 => "000011011000",
    3375 => "000011011001",
    3376 => "000011011010",
    3377 => "000011011100",
    3378 => "000011011101",
    3379 => "000011011111",
    3380 => "000011100000",
    3381 => "000011100010",
    3382 => "000011100011",
    3383 => "000011100100",
    3384 => "000011100110",
    3385 => "000011100111",
    3386 => "000011101001",
    3387 => "000011101010",
    3388 => "000011101100",
    3389 => "000011101101",
    3390 => "000011101111",
    3391 => "000011110000",
    3392 => "000011110010",
    3393 => "000011110011",
    3394 => "000011110101",
    3395 => "000011110110",
    3396 => "000011111000",
    3397 => "000011111001",
    3398 => "000011111011",
    3399 => "000011111100",
    3400 => "000011111110",
    3401 => "000011111111",
    3402 => "000100000001",
    3403 => "000100000010",
    3404 => "000100000100",
    3405 => "000100000101",
    3406 => "000100000111",
    3407 => "000100001000",
    3408 => "000100001010",
    3409 => "000100001011",
    3410 => "000100001101",
    3411 => "000100001110",
    3412 => "000100010000",
    3413 => "000100010010",
    3414 => "000100010011",
    3415 => "000100010101",
    3416 => "000100010110",
    3417 => "000100011000",
    3418 => "000100011001",
    3419 => "000100011011",
    3420 => "000100011101",
    3421 => "000100011110",
    3422 => "000100100000",
    3423 => "000100100001",
    3424 => "000100100011",
    3425 => "000100100101",
    3426 => "000100100110",
    3427 => "000100101000",
    3428 => "000100101010",
    3429 => "000100101011",
    3430 => "000100101101",
    3431 => "000100101110",
    3432 => "000100110000",
    3433 => "000100110010",
    3434 => "000100110011",
    3435 => "000100110101",
    3436 => "000100110111",
    3437 => "000100111000",
    3438 => "000100111010",
    3439 => "000100111100",
    3440 => "000100111101",
    3441 => "000100111111",
    3442 => "000101000001",
    3443 => "000101000010",
    3444 => "000101000100",
    3445 => "000101000110",
    3446 => "000101001000",
    3447 => "000101001001",
    3448 => "000101001011",
    3449 => "000101001101",
    3450 => "000101001110",
    3451 => "000101010000",
    3452 => "000101010010",
    3453 => "000101010100",
    3454 => "000101010101",
    3455 => "000101010111",
    3456 => "000101011001",
    3457 => "000101011011",
    3458 => "000101011100",
    3459 => "000101011110",
    3460 => "000101100000",
    3461 => "000101100010",
    3462 => "000101100011",
    3463 => "000101100101",
    3464 => "000101100111",
    3465 => "000101101001",
    3466 => "000101101010",
    3467 => "000101101100",
    3468 => "000101101110",
    3469 => "000101110000",
    3470 => "000101110010",
    3471 => "000101110011",
    3472 => "000101110101",
    3473 => "000101110111",
    3474 => "000101111001",
    3475 => "000101111011",
    3476 => "000101111101",
    3477 => "000101111110",
    3478 => "000110000000",
    3479 => "000110000010",
    3480 => "000110000100",
    3481 => "000110000110",
    3482 => "000110001000",
    3483 => "000110001001",
    3484 => "000110001011",
    3485 => "000110001101",
    3486 => "000110001111",
    3487 => "000110010001",
    3488 => "000110010011",
    3489 => "000110010101",
    3490 => "000110010110",
    3491 => "000110011000",
    3492 => "000110011010",
    3493 => "000110011100",
    3494 => "000110011110",
    3495 => "000110100000",
    3496 => "000110100010",
    3497 => "000110100100",
    3498 => "000110100110",
    3499 => "000110100111",
    3500 => "000110101001",
    3501 => "000110101011",
    3502 => "000110101101",
    3503 => "000110101111",
    3504 => "000110110001",
    3505 => "000110110011",
    3506 => "000110110101",
    3507 => "000110110111",
    3508 => "000110111001",
    3509 => "000110111011",
    3510 => "000110111101",
    3511 => "000110111111",
    3512 => "000111000001",
    3513 => "000111000011",
    3514 => "000111000101",
    3515 => "000111000111",
    3516 => "000111001001",
    3517 => "000111001011",
    3518 => "000111001101",
    3519 => "000111001111",
    3520 => "000111010001",
    3521 => "000111010011",
    3522 => "000111010100",
    3523 => "000111010111",
    3524 => "000111011001",
    3525 => "000111011011",
    3526 => "000111011101",
    3527 => "000111011111",
    3528 => "000111100001",
    3529 => "000111100011",
    3530 => "000111100101",
    3531 => "000111100111",
    3532 => "000111101001",
    3533 => "000111101011",
    3534 => "000111101101",
    3535 => "000111101111",
    3536 => "000111110001",
    3537 => "000111110011",
    3538 => "000111110101",
    3539 => "000111110111",
    3540 => "000111111001",
    3541 => "000111111011",
    3542 => "000111111101",
    3543 => "000111111111",
    3544 => "001000000001",
    3545 => "001000000011",
    3546 => "001000000110",
    3547 => "001000001000",
    3548 => "001000001010",
    3549 => "001000001100",
    3550 => "001000001110",
    3551 => "001000010000",
    3552 => "001000010010",
    3553 => "001000010100",
    3554 => "001000010110",
    3555 => "001000011000",
    3556 => "001000011011",
    3557 => "001000011101",
    3558 => "001000011111",
    3559 => "001000100001",
    3560 => "001000100011",
    3561 => "001000100101",
    3562 => "001000100111",
    3563 => "001000101010",
    3564 => "001000101100",
    3565 => "001000101110",
    3566 => "001000110000",
    3567 => "001000110010",
    3568 => "001000110100",
    3569 => "001000110111",
    3570 => "001000111001",
    3571 => "001000111011",
    3572 => "001000111101",
    3573 => "001000111111",
    3574 => "001001000001",
    3575 => "001001000100",
    3576 => "001001000110",
    3577 => "001001001000",
    3578 => "001001001010",
    3579 => "001001001100",
    3580 => "001001001111",
    3581 => "001001010001",
    3582 => "001001010011",
    3583 => "001001010101",
    3584 => "001001010111",
    3585 => "001001011010",
    3586 => "001001011100",
    3587 => "001001011110",
    3588 => "001001100000",
    3589 => "001001100011",
    3590 => "001001100101",
    3591 => "001001100111",
    3592 => "001001101001",
    3593 => "001001101100",
    3594 => "001001101110",
    3595 => "001001110000",
    3596 => "001001110010",
    3597 => "001001110101",
    3598 => "001001110111",
    3599 => "001001111001",
    3600 => "001001111011",
    3601 => "001001111110",
    3602 => "001010000000",
    3603 => "001010000010",
    3604 => "001010000101",
    3605 => "001010000111",
    3606 => "001010001001",
    3607 => "001010001011",
    3608 => "001010001110",
    3609 => "001010010000",
    3610 => "001010010010",
    3611 => "001010010101",
    3612 => "001010010111",
    3613 => "001010011001",
    3614 => "001010011100",
    3615 => "001010011110",
    3616 => "001010100000",
    3617 => "001010100011",
    3618 => "001010100101",
    3619 => "001010100111",
    3620 => "001010101010",
    3621 => "001010101100",
    3622 => "001010101110",
    3623 => "001010110001",
    3624 => "001010110011",
    3625 => "001010110101",
    3626 => "001010111000",
    3627 => "001010111010",
    3628 => "001010111100",
    3629 => "001010111111",
    3630 => "001011000001",
    3631 => "001011000011",
    3632 => "001011000110",
    3633 => "001011001000",
    3634 => "001011001011",
    3635 => "001011001101",
    3636 => "001011001111",
    3637 => "001011010010",
    3638 => "001011010100",
    3639 => "001011010111",
    3640 => "001011011001",
    3641 => "001011011011",
    3642 => "001011011110",
    3643 => "001011100000",
    3644 => "001011100011",
    3645 => "001011100101",
    3646 => "001011100111",
    3647 => "001011101010",
    3648 => "001011101100",
    3649 => "001011101111",
    3650 => "001011110001",
    3651 => "001011110100",
    3652 => "001011110110",
    3653 => "001011111000",
    3654 => "001011111011",
    3655 => "001011111101",
    3656 => "001100000000",
    3657 => "001100000010",
    3658 => "001100000101",
    3659 => "001100000111",
    3660 => "001100001010",
    3661 => "001100001100",
    3662 => "001100001111",
    3663 => "001100010001",
    3664 => "001100010100",
    3665 => "001100010110",
    3666 => "001100011000",
    3667 => "001100011011",
    3668 => "001100011101",
    3669 => "001100100000",
    3670 => "001100100010",
    3671 => "001100100101",
    3672 => "001100100111",
    3673 => "001100101010",
    3674 => "001100101100",
    3675 => "001100101111",
    3676 => "001100110001",
    3677 => "001100110100",
    3678 => "001100110110",
    3679 => "001100111001",
    3680 => "001100111011",
    3681 => "001100111110",
    3682 => "001101000001",
    3683 => "001101000011",
    3684 => "001101000110",
    3685 => "001101001000",
    3686 => "001101001011",
    3687 => "001101001101",
    3688 => "001101010000",
    3689 => "001101010010",
    3690 => "001101010101",
    3691 => "001101010111",
    3692 => "001101011010",
    3693 => "001101011101",
    3694 => "001101011111",
    3695 => "001101100010",
    3696 => "001101100100",
    3697 => "001101100111",
    3698 => "001101101001",
    3699 => "001101101100",
    3700 => "001101101111",
    3701 => "001101110001",
    3702 => "001101110100",
    3703 => "001101110110",
    3704 => "001101111001",
    3705 => "001101111011",
    3706 => "001101111110",
    3707 => "001110000001",
    3708 => "001110000011",
    3709 => "001110000110",
    3710 => "001110001000",
    3711 => "001110001011",
    3712 => "001110001110",
    3713 => "001110010000",
    3714 => "001110010011",
    3715 => "001110010101",
    3716 => "001110011000",
    3717 => "001110011011",
    3718 => "001110011101",
    3719 => "001110100000",
    3720 => "001110100011",
    3721 => "001110100101",
    3722 => "001110101000",
    3723 => "001110101011",
    3724 => "001110101101",
    3725 => "001110110000",
    3726 => "001110110010",
    3727 => "001110110101",
    3728 => "001110111000",
    3729 => "001110111010",
    3730 => "001110111101",
    3731 => "001111000000",
    3732 => "001111000010",
    3733 => "001111000101",
    3734 => "001111001000",
    3735 => "001111001010",
    3736 => "001111001101",
    3737 => "001111010000",
    3738 => "001111010010",
    3739 => "001111010101",
    3740 => "001111011000",
    3741 => "001111011010",
    3742 => "001111011101",
    3743 => "001111100000",
    3744 => "001111100011",
    3745 => "001111100101",
    3746 => "001111101000",
    3747 => "001111101011",
    3748 => "001111101101",
    3749 => "001111110000",
    3750 => "001111110011",
    3751 => "001111110101",
    3752 => "001111111000",
    3753 => "001111111011",
    3754 => "001111111110",
    3755 => "010000000000",
    3756 => "010000000011",
    3757 => "010000000110",
    3758 => "010000001000",
    3759 => "010000001011",
    3760 => "010000001110",
    3761 => "010000010001",
    3762 => "010000010011",
    3763 => "010000010110",
    3764 => "010000011001",
    3765 => "010000011100",
    3766 => "010000011110",
    3767 => "010000100001",
    3768 => "010000100100",
    3769 => "010000100111",
    3770 => "010000101001",
    3771 => "010000101100",
    3772 => "010000101111",
    3773 => "010000110010",
    3774 => "010000110100",
    3775 => "010000110111",
    3776 => "010000111010",
    3777 => "010000111101",
    3778 => "010001000000",
    3779 => "010001000010",
    3780 => "010001000101",
    3781 => "010001001000",
    3782 => "010001001011",
    3783 => "010001001101",
    3784 => "010001010000",
    3785 => "010001010011",
    3786 => "010001010110",
    3787 => "010001011001",
    3788 => "010001011011",
    3789 => "010001011110",
    3790 => "010001100001",
    3791 => "010001100100",
    3792 => "010001100111",
    3793 => "010001101001",
    3794 => "010001101100",
    3795 => "010001101111",
    3796 => "010001110010",
    3797 => "010001110101",
    3798 => "010001110111",
    3799 => "010001111010",
    3800 => "010001111101",
    3801 => "010010000000",
    3802 => "010010000011",
    3803 => "010010000110",
    3804 => "010010001000",
    3805 => "010010001011",
    3806 => "010010001110",
    3807 => "010010010001",
    3808 => "010010010100",
    3809 => "010010010111",
    3810 => "010010011001",
    3811 => "010010011100",
    3812 => "010010011111",
    3813 => "010010100010",
    3814 => "010010100101",
    3815 => "010010101000",
    3816 => "010010101010",
    3817 => "010010101101",
    3818 => "010010110000",
    3819 => "010010110011",
    3820 => "010010110110",
    3821 => "010010111001",
    3822 => "010010111100",
    3823 => "010010111111",
    3824 => "010011000001",
    3825 => "010011000100",
    3826 => "010011000111",
    3827 => "010011001010",
    3828 => "010011001101",
    3829 => "010011010000",
    3830 => "010011010011",
    3831 => "010011010110",
    3832 => "010011011000",
    3833 => "010011011011",
    3834 => "010011011110",
    3835 => "010011100001",
    3836 => "010011100100",
    3837 => "010011100111",
    3838 => "010011101010",
    3839 => "010011101101",
    3840 => "010011110000",
    3841 => "010011110010",
    3842 => "010011110101",
    3843 => "010011111000",
    3844 => "010011111011",
    3845 => "010011111110",
    3846 => "010100000001",
    3847 => "010100000100",
    3848 => "010100000111",
    3849 => "010100001010",
    3850 => "010100001101",
    3851 => "010100010000",
    3852 => "010100010011",
    3853 => "010100010101",
    3854 => "010100011000",
    3855 => "010100011011",
    3856 => "010100011110",
    3857 => "010100100001",
    3858 => "010100100100",
    3859 => "010100100111",
    3860 => "010100101010",
    3861 => "010100101101",
    3862 => "010100110000",
    3863 => "010100110011",
    3864 => "010100110110",
    3865 => "010100111001",
    3866 => "010100111100",
    3867 => "010100111111",
    3868 => "010101000010",
    3869 => "010101000100",
    3870 => "010101000111",
    3871 => "010101001010",
    3872 => "010101001101",
    3873 => "010101010000",
    3874 => "010101010011",
    3875 => "010101010110",
    3876 => "010101011001",
    3877 => "010101011100",
    3878 => "010101011111",
    3879 => "010101100010",
    3880 => "010101100101",
    3881 => "010101101000",
    3882 => "010101101011",
    3883 => "010101101110",
    3884 => "010101110001",
    3885 => "010101110100",
    3886 => "010101110111",
    3887 => "010101111010",
    3888 => "010101111101",
    3889 => "010110000000",
    3890 => "010110000011",
    3891 => "010110000110",
    3892 => "010110001001",
    3893 => "010110001100",
    3894 => "010110001111",
    3895 => "010110010010",
    3896 => "010110010101",
    3897 => "010110011000",
    3898 => "010110011011",
    3899 => "010110011110",
    3900 => "010110100001",
    3901 => "010110100100",
    3902 => "010110100111",
    3903 => "010110101010",
    3904 => "010110101101",
    3905 => "010110110000",
    3906 => "010110110011",
    3907 => "010110110110",
    3908 => "010110111001",
    3909 => "010110111100",
    3910 => "010110111111",
    3911 => "010111000010",
    3912 => "010111000101",
    3913 => "010111001000",
    3914 => "010111001011",
    3915 => "010111001110",
    3916 => "010111010001",
    3917 => "010111010100",
    3918 => "010111010111",
    3919 => "010111011010",
    3920 => "010111011101",
    3921 => "010111100000",
    3922 => "010111100011",
    3923 => "010111100110",
    3924 => "010111101001",
    3925 => "010111101100",
    3926 => "010111101111",
    3927 => "010111110010",
    3928 => "010111110101",
    3929 => "010111111000",
    3930 => "010111111011",
    3931 => "010111111110",
    3932 => "011000000001",
    3933 => "011000000100",
    3934 => "011000000111",
    3935 => "011000001011",
    3936 => "011000001110",
    3937 => "011000010001",
    3938 => "011000010100",
    3939 => "011000010111",
    3940 => "011000011010",
    3941 => "011000011101",
    3942 => "011000100000",
    3943 => "011000100011",
    3944 => "011000100110",
    3945 => "011000101001",
    3946 => "011000101100",
    3947 => "011000101111",
    3948 => "011000110010",
    3949 => "011000110101",
    3950 => "011000111000",
    3951 => "011000111011",
    3952 => "011000111110",
    3953 => "011001000010",
    3954 => "011001000101",
    3955 => "011001001000",
    3956 => "011001001011",
    3957 => "011001001110",
    3958 => "011001010001",
    3959 => "011001010100",
    3960 => "011001010111",
    3961 => "011001011010",
    3962 => "011001011101",
    3963 => "011001100000",
    3964 => "011001100011",
    3965 => "011001100110",
    3966 => "011001101001",
    3967 => "011001101101",
    3968 => "011001110000",
    3969 => "011001110011",
    3970 => "011001110110",
    3971 => "011001111001",
    3972 => "011001111100",
    3973 => "011001111111",
    3974 => "011010000010",
    3975 => "011010000101",
    3976 => "011010001000",
    3977 => "011010001011",
    3978 => "011010001110",
    3979 => "011010010010",
    3980 => "011010010101",
    3981 => "011010011000",
    3982 => "011010011011",
    3983 => "011010011110",
    3984 => "011010100001",
    3985 => "011010100100",
    3986 => "011010100111",
    3987 => "011010101010",
    3988 => "011010101101",
    3989 => "011010110000",
    3990 => "011010110100",
    3991 => "011010110111",
    3992 => "011010111010",
    3993 => "011010111101",
    3994 => "011011000000",
    3995 => "011011000011",
    3996 => "011011000110",
    3997 => "011011001001",
    3998 => "011011001100",
    3999 => "011011010000",
    4000 => "011011010011",
    4001 => "011011010110",
    4002 => "011011011001",
    4003 => "011011011100",
    4004 => "011011011111",
    4005 => "011011100010",
    4006 => "011011100101",
    4007 => "011011101000",
    4008 => "011011101011",
    4009 => "011011101111",
    4010 => "011011110010",
    4011 => "011011110101",
    4012 => "011011111000",
    4013 => "011011111011",
    4014 => "011011111110",
    4015 => "011100000001",
    4016 => "011100000100",
    4017 => "011100001000",
    4018 => "011100001011",
    4019 => "011100001110",
    4020 => "011100010001",
    4021 => "011100010100",
    4022 => "011100010111",
    4023 => "011100011010",
    4024 => "011100011101",
    4025 => "011100100000",
    4026 => "011100100100",
    4027 => "011100100111",
    4028 => "011100101010",
    4029 => "011100101101",
    4030 => "011100110000",
    4031 => "011100110011",
    4032 => "011100110110",
    4033 => "011100111001",
    4034 => "011100111101",
    4035 => "011101000000",
    4036 => "011101000011",
    4037 => "011101000110",
    4038 => "011101001001",
    4039 => "011101001100",
    4040 => "011101001111",
    4041 => "011101010010",
    4042 => "011101010110",
    4043 => "011101011001",
    4044 => "011101011100",
    4045 => "011101011111",
    4046 => "011101100010",
    4047 => "011101100101",
    4048 => "011101101000",
    4049 => "011101101100",
    4050 => "011101101111",
    4051 => "011101110010",
    4052 => "011101110101",
    4053 => "011101111000",
    4054 => "011101111011",
    4055 => "011101111110",
    4056 => "011110000001",
    4057 => "011110000101",
    4058 => "011110001000",
    4059 => "011110001011",
    4060 => "011110001110",
    4061 => "011110010001",
    4062 => "011110010100",
    4063 => "011110010111",
    4064 => "011110011011",
    4065 => "011110011110",
    4066 => "011110100001",
    4067 => "011110100100",
    4068 => "011110100111",
    4069 => "011110101010",
    4070 => "011110101101",
    4071 => "011110110001",
    4072 => "011110110100",
    4073 => "011110110111",
    4074 => "011110111010",
    4075 => "011110111101",
    4076 => "011111000000",
    4077 => "011111000011",
    4078 => "011111000110",
    4079 => "011111001010",
    4080 => "011111001101",
    4081 => "011111010000",
    4082 => "011111010011",
    4083 => "011111010110",
    4084 => "011111011001",
    4085 => "011111011100",
    4086 => "011111100000",
    4087 => "011111100011",
    4088 => "011111100110",
    4089 => "011111101001",
    4090 => "011111101100",
    4091 => "011111101111",
    4092 => "011111110010",
    4093 => "011111110110",
    4094 => "011111111001",
    4095 => "011111111001");
begin
 process (address)
 begin
  case address is
     when "000000000000" => data <= sine_rom(0);
     when "000000000001" => data <= sine_rom(1);
     when "000000000010" => data <= sine_rom(2);
     when "000000000011" => data <= sine_rom(3);
     when "000000000100" => data <= sine_rom(4);
     when "000000000101" => data <= sine_rom(5);
     when "000000000110" => data <= sine_rom(6);
     when "000000000111" => data <= sine_rom(7);
     when "000000001000" => data <= sine_rom(8);
     when "000000001001" => data <= sine_rom(9);
     when "000000001010" => data <= sine_rom(10);
     when "000000001011" => data <= sine_rom(11);
     when "000000001100" => data <= sine_rom(12);
     when "000000001101" => data <= sine_rom(13);
     when "000000001110" => data <= sine_rom(14);
     when "000000001111" => data <= sine_rom(15);
     when "000000010000" => data <= sine_rom(16);
     when "000000010001" => data <= sine_rom(17);
     when "000000010010" => data <= sine_rom(18);
     when "000000010011" => data <= sine_rom(19);
     when "000000010100" => data <= sine_rom(20);
     when "000000010101" => data <= sine_rom(21);
     when "000000010110" => data <= sine_rom(22);
     when "000000010111" => data <= sine_rom(23);
     when "000000011000" => data <= sine_rom(24);
     when "000000011001" => data <= sine_rom(25);
     when "000000011010" => data <= sine_rom(26);
     when "000000011011" => data <= sine_rom(27);
     when "000000011100" => data <= sine_rom(28);
     when "000000011101" => data <= sine_rom(29);
     when "000000011110" => data <= sine_rom(30);
     when "000000011111" => data <= sine_rom(31);
     when "000000100000" => data <= sine_rom(32);
     when "000000100001" => data <= sine_rom(33);
     when "000000100010" => data <= sine_rom(34);
     when "000000100011" => data <= sine_rom(35);
     when "000000100100" => data <= sine_rom(36);
     when "000000100101" => data <= sine_rom(37);
     when "000000100110" => data <= sine_rom(38);
     when "000000100111" => data <= sine_rom(39);
     when "000000101000" => data <= sine_rom(40);
     when "000000101001" => data <= sine_rom(41);
     when "000000101010" => data <= sine_rom(42);
     when "000000101011" => data <= sine_rom(43);
     when "000000101100" => data <= sine_rom(44);
     when "000000101101" => data <= sine_rom(45);
     when "000000101110" => data <= sine_rom(46);
     when "000000101111" => data <= sine_rom(47);
     when "000000110000" => data <= sine_rom(48);
     when "000000110001" => data <= sine_rom(49);
     when "000000110010" => data <= sine_rom(50);
     when "000000110011" => data <= sine_rom(51);
     when "000000110100" => data <= sine_rom(52);
     when "000000110101" => data <= sine_rom(53);
     when "000000110110" => data <= sine_rom(54);
     when "000000110111" => data <= sine_rom(55);
     when "000000111000" => data <= sine_rom(56);
     when "000000111001" => data <= sine_rom(57);
     when "000000111010" => data <= sine_rom(58);
     when "000000111011" => data <= sine_rom(59);
     when "000000111100" => data <= sine_rom(60);
     when "000000111101" => data <= sine_rom(61);
     when "000000111110" => data <= sine_rom(62);
     when "000000111111" => data <= sine_rom(63);
     when "000001000000" => data <= sine_rom(64);
     when "000001000001" => data <= sine_rom(65);
     when "000001000010" => data <= sine_rom(66);
     when "000001000011" => data <= sine_rom(67);
     when "000001000100" => data <= sine_rom(68);
     when "000001000101" => data <= sine_rom(69);
     when "000001000110" => data <= sine_rom(70);
     when "000001000111" => data <= sine_rom(71);
     when "000001001000" => data <= sine_rom(72);
     when "000001001001" => data <= sine_rom(73);
     when "000001001010" => data <= sine_rom(74);
     when "000001001011" => data <= sine_rom(75);
     when "000001001100" => data <= sine_rom(76);
     when "000001001101" => data <= sine_rom(77);
     when "000001001110" => data <= sine_rom(78);
     when "000001001111" => data <= sine_rom(79);
     when "000001010000" => data <= sine_rom(80);
     when "000001010001" => data <= sine_rom(81);
     when "000001010010" => data <= sine_rom(82);
     when "000001010011" => data <= sine_rom(83);
     when "000001010100" => data <= sine_rom(84);
     when "000001010101" => data <= sine_rom(85);
     when "000001010110" => data <= sine_rom(86);
     when "000001010111" => data <= sine_rom(87);
     when "000001011000" => data <= sine_rom(88);
     when "000001011001" => data <= sine_rom(89);
     when "000001011010" => data <= sine_rom(90);
     when "000001011011" => data <= sine_rom(91);
     when "000001011100" => data <= sine_rom(92);
     when "000001011101" => data <= sine_rom(93);
     when "000001011110" => data <= sine_rom(94);
     when "000001011111" => data <= sine_rom(95);
     when "000001100000" => data <= sine_rom(96);
     when "000001100001" => data <= sine_rom(97);
     when "000001100010" => data <= sine_rom(98);
     when "000001100011" => data <= sine_rom(99);
     when "000001100100" => data <= sine_rom(100);
     when "000001100101" => data <= sine_rom(101);
     when "000001100110" => data <= sine_rom(102);
     when "000001100111" => data <= sine_rom(103);
     when "000001101000" => data <= sine_rom(104);
     when "000001101001" => data <= sine_rom(105);
     when "000001101010" => data <= sine_rom(106);
     when "000001101011" => data <= sine_rom(107);
     when "000001101100" => data <= sine_rom(108);
     when "000001101101" => data <= sine_rom(109);
     when "000001101110" => data <= sine_rom(110);
     when "000001101111" => data <= sine_rom(111);
     when "000001110000" => data <= sine_rom(112);
     when "000001110001" => data <= sine_rom(113);
     when "000001110010" => data <= sine_rom(114);
     when "000001110011" => data <= sine_rom(115);
     when "000001110100" => data <= sine_rom(116);
     when "000001110101" => data <= sine_rom(117);
     when "000001110110" => data <= sine_rom(118);
     when "000001110111" => data <= sine_rom(119);
     when "000001111000" => data <= sine_rom(120);
     when "000001111001" => data <= sine_rom(121);
     when "000001111010" => data <= sine_rom(122);
     when "000001111011" => data <= sine_rom(123);
     when "000001111100" => data <= sine_rom(124);
     when "000001111101" => data <= sine_rom(125);
     when "000001111110" => data <= sine_rom(126);
     when "000001111111" => data <= sine_rom(127);
     when "000010000000" => data <= sine_rom(128);
     when "000010000001" => data <= sine_rom(129);
     when "000010000010" => data <= sine_rom(130);
     when "000010000011" => data <= sine_rom(131);
     when "000010000100" => data <= sine_rom(132);
     when "000010000101" => data <= sine_rom(133);
     when "000010000110" => data <= sine_rom(134);
     when "000010000111" => data <= sine_rom(135);
     when "000010001000" => data <= sine_rom(136);
     when "000010001001" => data <= sine_rom(137);
     when "000010001010" => data <= sine_rom(138);
     when "000010001011" => data <= sine_rom(139);
     when "000010001100" => data <= sine_rom(140);
     when "000010001101" => data <= sine_rom(141);
     when "000010001110" => data <= sine_rom(142);
     when "000010001111" => data <= sine_rom(143);
     when "000010010000" => data <= sine_rom(144);
     when "000010010001" => data <= sine_rom(145);
     when "000010010010" => data <= sine_rom(146);
     when "000010010011" => data <= sine_rom(147);
     when "000010010100" => data <= sine_rom(148);
     when "000010010101" => data <= sine_rom(149);
     when "000010010110" => data <= sine_rom(150);
     when "000010010111" => data <= sine_rom(151);
     when "000010011000" => data <= sine_rom(152);
     when "000010011001" => data <= sine_rom(153);
     when "000010011010" => data <= sine_rom(154);
     when "000010011011" => data <= sine_rom(155);
     when "000010011100" => data <= sine_rom(156);
     when "000010011101" => data <= sine_rom(157);
     when "000010011110" => data <= sine_rom(158);
     when "000010011111" => data <= sine_rom(159);
     when "000010100000" => data <= sine_rom(160);
     when "000010100001" => data <= sine_rom(161);
     when "000010100010" => data <= sine_rom(162);
     when "000010100011" => data <= sine_rom(163);
     when "000010100100" => data <= sine_rom(164);
     when "000010100101" => data <= sine_rom(165);
     when "000010100110" => data <= sine_rom(166);
     when "000010100111" => data <= sine_rom(167);
     when "000010101000" => data <= sine_rom(168);
     when "000010101001" => data <= sine_rom(169);
     when "000010101010" => data <= sine_rom(170);
     when "000010101011" => data <= sine_rom(171);
     when "000010101100" => data <= sine_rom(172);
     when "000010101101" => data <= sine_rom(173);
     when "000010101110" => data <= sine_rom(174);
     when "000010101111" => data <= sine_rom(175);
     when "000010110000" => data <= sine_rom(176);
     when "000010110001" => data <= sine_rom(177);
     when "000010110010" => data <= sine_rom(178);
     when "000010110011" => data <= sine_rom(179);
     when "000010110100" => data <= sine_rom(180);
     when "000010110101" => data <= sine_rom(181);
     when "000010110110" => data <= sine_rom(182);
     when "000010110111" => data <= sine_rom(183);
     when "000010111000" => data <= sine_rom(184);
     when "000010111001" => data <= sine_rom(185);
     when "000010111010" => data <= sine_rom(186);
     when "000010111011" => data <= sine_rom(187);
     when "000010111100" => data <= sine_rom(188);
     when "000010111101" => data <= sine_rom(189);
     when "000010111110" => data <= sine_rom(190);
     when "000010111111" => data <= sine_rom(191);
     when "000011000000" => data <= sine_rom(192);
     when "000011000001" => data <= sine_rom(193);
     when "000011000010" => data <= sine_rom(194);
     when "000011000011" => data <= sine_rom(195);
     when "000011000100" => data <= sine_rom(196);
     when "000011000101" => data <= sine_rom(197);
     when "000011000110" => data <= sine_rom(198);
     when "000011000111" => data <= sine_rom(199);
     when "000011001000" => data <= sine_rom(200);
     when "000011001001" => data <= sine_rom(201);
     when "000011001010" => data <= sine_rom(202);
     when "000011001011" => data <= sine_rom(203);
     when "000011001100" => data <= sine_rom(204);
     when "000011001101" => data <= sine_rom(205);
     when "000011001110" => data <= sine_rom(206);
     when "000011001111" => data <= sine_rom(207);
     when "000011010000" => data <= sine_rom(208);
     when "000011010001" => data <= sine_rom(209);
     when "000011010010" => data <= sine_rom(210);
     when "000011010011" => data <= sine_rom(211);
     when "000011010100" => data <= sine_rom(212);
     when "000011010101" => data <= sine_rom(213);
     when "000011010110" => data <= sine_rom(214);
     when "000011010111" => data <= sine_rom(215);
     when "000011011000" => data <= sine_rom(216);
     when "000011011001" => data <= sine_rom(217);
     when "000011011010" => data <= sine_rom(218);
     when "000011011011" => data <= sine_rom(219);
     when "000011011100" => data <= sine_rom(220);
     when "000011011101" => data <= sine_rom(221);
     when "000011011110" => data <= sine_rom(222);
     when "000011011111" => data <= sine_rom(223);
     when "000011100000" => data <= sine_rom(224);
     when "000011100001" => data <= sine_rom(225);
     when "000011100010" => data <= sine_rom(226);
     when "000011100011" => data <= sine_rom(227);
     when "000011100100" => data <= sine_rom(228);
     when "000011100101" => data <= sine_rom(229);
     when "000011100110" => data <= sine_rom(230);
     when "000011100111" => data <= sine_rom(231);
     when "000011101000" => data <= sine_rom(232);
     when "000011101001" => data <= sine_rom(233);
     when "000011101010" => data <= sine_rom(234);
     when "000011101011" => data <= sine_rom(235);
     when "000011101100" => data <= sine_rom(236);
     when "000011101101" => data <= sine_rom(237);
     when "000011101110" => data <= sine_rom(238);
     when "000011101111" => data <= sine_rom(239);
     when "000011110000" => data <= sine_rom(240);
     when "000011110001" => data <= sine_rom(241);
     when "000011110010" => data <= sine_rom(242);
     when "000011110011" => data <= sine_rom(243);
     when "000011110100" => data <= sine_rom(244);
     when "000011110101" => data <= sine_rom(245);
     when "000011110110" => data <= sine_rom(246);
     when "000011110111" => data <= sine_rom(247);
     when "000011111000" => data <= sine_rom(248);
     when "000011111001" => data <= sine_rom(249);
     when "000011111010" => data <= sine_rom(250);
     when "000011111011" => data <= sine_rom(251);
     when "000011111100" => data <= sine_rom(252);
     when "000011111101" => data <= sine_rom(253);
     when "000011111110" => data <= sine_rom(254);
     when "000011111111" => data <= sine_rom(255);
     when "000100000000" => data <= sine_rom(256);
     when "000100000001" => data <= sine_rom(257);
     when "000100000010" => data <= sine_rom(258);
     when "000100000011" => data <= sine_rom(259);
     when "000100000100" => data <= sine_rom(260);
     when "000100000101" => data <= sine_rom(261);
     when "000100000110" => data <= sine_rom(262);
     when "000100000111" => data <= sine_rom(263);
     when "000100001000" => data <= sine_rom(264);
     when "000100001001" => data <= sine_rom(265);
     when "000100001010" => data <= sine_rom(266);
     when "000100001011" => data <= sine_rom(267);
     when "000100001100" => data <= sine_rom(268);
     when "000100001101" => data <= sine_rom(269);
     when "000100001110" => data <= sine_rom(270);
     when "000100001111" => data <= sine_rom(271);
     when "000100010000" => data <= sine_rom(272);
     when "000100010001" => data <= sine_rom(273);
     when "000100010010" => data <= sine_rom(274);
     when "000100010011" => data <= sine_rom(275);
     when "000100010100" => data <= sine_rom(276);
     when "000100010101" => data <= sine_rom(277);
     when "000100010110" => data <= sine_rom(278);
     when "000100010111" => data <= sine_rom(279);
     when "000100011000" => data <= sine_rom(280);
     when "000100011001" => data <= sine_rom(281);
     when "000100011010" => data <= sine_rom(282);
     when "000100011011" => data <= sine_rom(283);
     when "000100011100" => data <= sine_rom(284);
     when "000100011101" => data <= sine_rom(285);
     when "000100011110" => data <= sine_rom(286);
     when "000100011111" => data <= sine_rom(287);
     when "000100100000" => data <= sine_rom(288);
     when "000100100001" => data <= sine_rom(289);
     when "000100100010" => data <= sine_rom(290);
     when "000100100011" => data <= sine_rom(291);
     when "000100100100" => data <= sine_rom(292);
     when "000100100101" => data <= sine_rom(293);
     when "000100100110" => data <= sine_rom(294);
     when "000100100111" => data <= sine_rom(295);
     when "000100101000" => data <= sine_rom(296);
     when "000100101001" => data <= sine_rom(297);
     when "000100101010" => data <= sine_rom(298);
     when "000100101011" => data <= sine_rom(299);
     when "000100101100" => data <= sine_rom(300);
     when "000100101101" => data <= sine_rom(301);
     when "000100101110" => data <= sine_rom(302);
     when "000100101111" => data <= sine_rom(303);
     when "000100110000" => data <= sine_rom(304);
     when "000100110001" => data <= sine_rom(305);
     when "000100110010" => data <= sine_rom(306);
     when "000100110011" => data <= sine_rom(307);
     when "000100110100" => data <= sine_rom(308);
     when "000100110101" => data <= sine_rom(309);
     when "000100110110" => data <= sine_rom(310);
     when "000100110111" => data <= sine_rom(311);
     when "000100111000" => data <= sine_rom(312);
     when "000100111001" => data <= sine_rom(313);
     when "000100111010" => data <= sine_rom(314);
     when "000100111011" => data <= sine_rom(315);
     when "000100111100" => data <= sine_rom(316);
     when "000100111101" => data <= sine_rom(317);
     when "000100111110" => data <= sine_rom(318);
     when "000100111111" => data <= sine_rom(319);
     when "000101000000" => data <= sine_rom(320);
     when "000101000001" => data <= sine_rom(321);
     when "000101000010" => data <= sine_rom(322);
     when "000101000011" => data <= sine_rom(323);
     when "000101000100" => data <= sine_rom(324);
     when "000101000101" => data <= sine_rom(325);
     when "000101000110" => data <= sine_rom(326);
     when "000101000111" => data <= sine_rom(327);
     when "000101001000" => data <= sine_rom(328);
     when "000101001001" => data <= sine_rom(329);
     when "000101001010" => data <= sine_rom(330);
     when "000101001011" => data <= sine_rom(331);
     when "000101001100" => data <= sine_rom(332);
     when "000101001101" => data <= sine_rom(333);
     when "000101001110" => data <= sine_rom(334);
     when "000101001111" => data <= sine_rom(335);
     when "000101010000" => data <= sine_rom(336);
     when "000101010001" => data <= sine_rom(337);
     when "000101010010" => data <= sine_rom(338);
     when "000101010011" => data <= sine_rom(339);
     when "000101010100" => data <= sine_rom(340);
     when "000101010101" => data <= sine_rom(341);
     when "000101010110" => data <= sine_rom(342);
     when "000101010111" => data <= sine_rom(343);
     when "000101011000" => data <= sine_rom(344);
     when "000101011001" => data <= sine_rom(345);
     when "000101011010" => data <= sine_rom(346);
     when "000101011011" => data <= sine_rom(347);
     when "000101011100" => data <= sine_rom(348);
     when "000101011101" => data <= sine_rom(349);
     when "000101011110" => data <= sine_rom(350);
     when "000101011111" => data <= sine_rom(351);
     when "000101100000" => data <= sine_rom(352);
     when "000101100001" => data <= sine_rom(353);
     when "000101100010" => data <= sine_rom(354);
     when "000101100011" => data <= sine_rom(355);
     when "000101100100" => data <= sine_rom(356);
     when "000101100101" => data <= sine_rom(357);
     when "000101100110" => data <= sine_rom(358);
     when "000101100111" => data <= sine_rom(359);
     when "000101101000" => data <= sine_rom(360);
     when "000101101001" => data <= sine_rom(361);
     when "000101101010" => data <= sine_rom(362);
     when "000101101011" => data <= sine_rom(363);
     when "000101101100" => data <= sine_rom(364);
     when "000101101101" => data <= sine_rom(365);
     when "000101101110" => data <= sine_rom(366);
     when "000101101111" => data <= sine_rom(367);
     when "000101110000" => data <= sine_rom(368);
     when "000101110001" => data <= sine_rom(369);
     when "000101110010" => data <= sine_rom(370);
     when "000101110011" => data <= sine_rom(371);
     when "000101110100" => data <= sine_rom(372);
     when "000101110101" => data <= sine_rom(373);
     when "000101110110" => data <= sine_rom(374);
     when "000101110111" => data <= sine_rom(375);
     when "000101111000" => data <= sine_rom(376);
     when "000101111001" => data <= sine_rom(377);
     when "000101111010" => data <= sine_rom(378);
     when "000101111011" => data <= sine_rom(379);
     when "000101111100" => data <= sine_rom(380);
     when "000101111101" => data <= sine_rom(381);
     when "000101111110" => data <= sine_rom(382);
     when "000101111111" => data <= sine_rom(383);
     when "000110000000" => data <= sine_rom(384);
     when "000110000001" => data <= sine_rom(385);
     when "000110000010" => data <= sine_rom(386);
     when "000110000011" => data <= sine_rom(387);
     when "000110000100" => data <= sine_rom(388);
     when "000110000101" => data <= sine_rom(389);
     when "000110000110" => data <= sine_rom(390);
     when "000110000111" => data <= sine_rom(391);
     when "000110001000" => data <= sine_rom(392);
     when "000110001001" => data <= sine_rom(393);
     when "000110001010" => data <= sine_rom(394);
     when "000110001011" => data <= sine_rom(395);
     when "000110001100" => data <= sine_rom(396);
     when "000110001101" => data <= sine_rom(397);
     when "000110001110" => data <= sine_rom(398);
     when "000110001111" => data <= sine_rom(399);
     when "000110010000" => data <= sine_rom(400);
     when "000110010001" => data <= sine_rom(401);
     when "000110010010" => data <= sine_rom(402);
     when "000110010011" => data <= sine_rom(403);
     when "000110010100" => data <= sine_rom(404);
     when "000110010101" => data <= sine_rom(405);
     when "000110010110" => data <= sine_rom(406);
     when "000110010111" => data <= sine_rom(407);
     when "000110011000" => data <= sine_rom(408);
     when "000110011001" => data <= sine_rom(409);
     when "000110011010" => data <= sine_rom(410);
     when "000110011011" => data <= sine_rom(411);
     when "000110011100" => data <= sine_rom(412);
     when "000110011101" => data <= sine_rom(413);
     when "000110011110" => data <= sine_rom(414);
     when "000110011111" => data <= sine_rom(415);
     when "000110100000" => data <= sine_rom(416);
     when "000110100001" => data <= sine_rom(417);
     when "000110100010" => data <= sine_rom(418);
     when "000110100011" => data <= sine_rom(419);
     when "000110100100" => data <= sine_rom(420);
     when "000110100101" => data <= sine_rom(421);
     when "000110100110" => data <= sine_rom(422);
     when "000110100111" => data <= sine_rom(423);
     when "000110101000" => data <= sine_rom(424);
     when "000110101001" => data <= sine_rom(425);
     when "000110101010" => data <= sine_rom(426);
     when "000110101011" => data <= sine_rom(427);
     when "000110101100" => data <= sine_rom(428);
     when "000110101101" => data <= sine_rom(429);
     when "000110101110" => data <= sine_rom(430);
     when "000110101111" => data <= sine_rom(431);
     when "000110110000" => data <= sine_rom(432);
     when "000110110001" => data <= sine_rom(433);
     when "000110110010" => data <= sine_rom(434);
     when "000110110011" => data <= sine_rom(435);
     when "000110110100" => data <= sine_rom(436);
     when "000110110101" => data <= sine_rom(437);
     when "000110110110" => data <= sine_rom(438);
     when "000110110111" => data <= sine_rom(439);
     when "000110111000" => data <= sine_rom(440);
     when "000110111001" => data <= sine_rom(441);
     when "000110111010" => data <= sine_rom(442);
     when "000110111011" => data <= sine_rom(443);
     when "000110111100" => data <= sine_rom(444);
     when "000110111101" => data <= sine_rom(445);
     when "000110111110" => data <= sine_rom(446);
     when "000110111111" => data <= sine_rom(447);
     when "000111000000" => data <= sine_rom(448);
     when "000111000001" => data <= sine_rom(449);
     when "000111000010" => data <= sine_rom(450);
     when "000111000011" => data <= sine_rom(451);
     when "000111000100" => data <= sine_rom(452);
     when "000111000101" => data <= sine_rom(453);
     when "000111000110" => data <= sine_rom(454);
     when "000111000111" => data <= sine_rom(455);
     when "000111001000" => data <= sine_rom(456);
     when "000111001001" => data <= sine_rom(457);
     when "000111001010" => data <= sine_rom(458);
     when "000111001011" => data <= sine_rom(459);
     when "000111001100" => data <= sine_rom(460);
     when "000111001101" => data <= sine_rom(461);
     when "000111001110" => data <= sine_rom(462);
     when "000111001111" => data <= sine_rom(463);
     when "000111010000" => data <= sine_rom(464);
     when "000111010001" => data <= sine_rom(465);
     when "000111010010" => data <= sine_rom(466);
     when "000111010011" => data <= sine_rom(467);
     when "000111010100" => data <= sine_rom(468);
     when "000111010101" => data <= sine_rom(469);
     when "000111010110" => data <= sine_rom(470);
     when "000111010111" => data <= sine_rom(471);
     when "000111011000" => data <= sine_rom(472);
     when "000111011001" => data <= sine_rom(473);
     when "000111011010" => data <= sine_rom(474);
     when "000111011011" => data <= sine_rom(475);
     when "000111011100" => data <= sine_rom(476);
     when "000111011101" => data <= sine_rom(477);
     when "000111011110" => data <= sine_rom(478);
     when "000111011111" => data <= sine_rom(479);
     when "000111100000" => data <= sine_rom(480);
     when "000111100001" => data <= sine_rom(481);
     when "000111100010" => data <= sine_rom(482);
     when "000111100011" => data <= sine_rom(483);
     when "000111100100" => data <= sine_rom(484);
     when "000111100101" => data <= sine_rom(485);
     when "000111100110" => data <= sine_rom(486);
     when "000111100111" => data <= sine_rom(487);
     when "000111101000" => data <= sine_rom(488);
     when "000111101001" => data <= sine_rom(489);
     when "000111101010" => data <= sine_rom(490);
     when "000111101011" => data <= sine_rom(491);
     when "000111101100" => data <= sine_rom(492);
     when "000111101101" => data <= sine_rom(493);
     when "000111101110" => data <= sine_rom(494);
     when "000111101111" => data <= sine_rom(495);
     when "000111110000" => data <= sine_rom(496);
     when "000111110001" => data <= sine_rom(497);
     when "000111110010" => data <= sine_rom(498);
     when "000111110011" => data <= sine_rom(499);
     when "000111110100" => data <= sine_rom(500);
     when "000111110101" => data <= sine_rom(501);
     when "000111110110" => data <= sine_rom(502);
     when "000111110111" => data <= sine_rom(503);
     when "000111111000" => data <= sine_rom(504);
     when "000111111001" => data <= sine_rom(505);
     when "000111111010" => data <= sine_rom(506);
     when "000111111011" => data <= sine_rom(507);
     when "000111111100" => data <= sine_rom(508);
     when "000111111101" => data <= sine_rom(509);
     when "000111111110" => data <= sine_rom(510);
     when "000111111111" => data <= sine_rom(511);
     when "001000000000" => data <= sine_rom(512);
     when "001000000001" => data <= sine_rom(513);
     when "001000000010" => data <= sine_rom(514);
     when "001000000011" => data <= sine_rom(515);
     when "001000000100" => data <= sine_rom(516);
     when "001000000101" => data <= sine_rom(517);
     when "001000000110" => data <= sine_rom(518);
     when "001000000111" => data <= sine_rom(519);
     when "001000001000" => data <= sine_rom(520);
     when "001000001001" => data <= sine_rom(521);
     when "001000001010" => data <= sine_rom(522);
     when "001000001011" => data <= sine_rom(523);
     when "001000001100" => data <= sine_rom(524);
     when "001000001101" => data <= sine_rom(525);
     when "001000001110" => data <= sine_rom(526);
     when "001000001111" => data <= sine_rom(527);
     when "001000010000" => data <= sine_rom(528);
     when "001000010001" => data <= sine_rom(529);
     when "001000010010" => data <= sine_rom(530);
     when "001000010011" => data <= sine_rom(531);
     when "001000010100" => data <= sine_rom(532);
     when "001000010101" => data <= sine_rom(533);
     when "001000010110" => data <= sine_rom(534);
     when "001000010111" => data <= sine_rom(535);
     when "001000011000" => data <= sine_rom(536);
     when "001000011001" => data <= sine_rom(537);
     when "001000011010" => data <= sine_rom(538);
     when "001000011011" => data <= sine_rom(539);
     when "001000011100" => data <= sine_rom(540);
     when "001000011101" => data <= sine_rom(541);
     when "001000011110" => data <= sine_rom(542);
     when "001000011111" => data <= sine_rom(543);
     when "001000100000" => data <= sine_rom(544);
     when "001000100001" => data <= sine_rom(545);
     when "001000100010" => data <= sine_rom(546);
     when "001000100011" => data <= sine_rom(547);
     when "001000100100" => data <= sine_rom(548);
     when "001000100101" => data <= sine_rom(549);
     when "001000100110" => data <= sine_rom(550);
     when "001000100111" => data <= sine_rom(551);
     when "001000101000" => data <= sine_rom(552);
     when "001000101001" => data <= sine_rom(553);
     when "001000101010" => data <= sine_rom(554);
     when "001000101011" => data <= sine_rom(555);
     when "001000101100" => data <= sine_rom(556);
     when "001000101101" => data <= sine_rom(557);
     when "001000101110" => data <= sine_rom(558);
     when "001000101111" => data <= sine_rom(559);
     when "001000110000" => data <= sine_rom(560);
     when "001000110001" => data <= sine_rom(561);
     when "001000110010" => data <= sine_rom(562);
     when "001000110011" => data <= sine_rom(563);
     when "001000110100" => data <= sine_rom(564);
     when "001000110101" => data <= sine_rom(565);
     when "001000110110" => data <= sine_rom(566);
     when "001000110111" => data <= sine_rom(567);
     when "001000111000" => data <= sine_rom(568);
     when "001000111001" => data <= sine_rom(569);
     when "001000111010" => data <= sine_rom(570);
     when "001000111011" => data <= sine_rom(571);
     when "001000111100" => data <= sine_rom(572);
     when "001000111101" => data <= sine_rom(573);
     when "001000111110" => data <= sine_rom(574);
     when "001000111111" => data <= sine_rom(575);
     when "001001000000" => data <= sine_rom(576);
     when "001001000001" => data <= sine_rom(577);
     when "001001000010" => data <= sine_rom(578);
     when "001001000011" => data <= sine_rom(579);
     when "001001000100" => data <= sine_rom(580);
     when "001001000101" => data <= sine_rom(581);
     when "001001000110" => data <= sine_rom(582);
     when "001001000111" => data <= sine_rom(583);
     when "001001001000" => data <= sine_rom(584);
     when "001001001001" => data <= sine_rom(585);
     when "001001001010" => data <= sine_rom(586);
     when "001001001011" => data <= sine_rom(587);
     when "001001001100" => data <= sine_rom(588);
     when "001001001101" => data <= sine_rom(589);
     when "001001001110" => data <= sine_rom(590);
     when "001001001111" => data <= sine_rom(591);
     when "001001010000" => data <= sine_rom(592);
     when "001001010001" => data <= sine_rom(593);
     when "001001010010" => data <= sine_rom(594);
     when "001001010011" => data <= sine_rom(595);
     when "001001010100" => data <= sine_rom(596);
     when "001001010101" => data <= sine_rom(597);
     when "001001010110" => data <= sine_rom(598);
     when "001001010111" => data <= sine_rom(599);
     when "001001011000" => data <= sine_rom(600);
     when "001001011001" => data <= sine_rom(601);
     when "001001011010" => data <= sine_rom(602);
     when "001001011011" => data <= sine_rom(603);
     when "001001011100" => data <= sine_rom(604);
     when "001001011101" => data <= sine_rom(605);
     when "001001011110" => data <= sine_rom(606);
     when "001001011111" => data <= sine_rom(607);
     when "001001100000" => data <= sine_rom(608);
     when "001001100001" => data <= sine_rom(609);
     when "001001100010" => data <= sine_rom(610);
     when "001001100011" => data <= sine_rom(611);
     when "001001100100" => data <= sine_rom(612);
     when "001001100101" => data <= sine_rom(613);
     when "001001100110" => data <= sine_rom(614);
     when "001001100111" => data <= sine_rom(615);
     when "001001101000" => data <= sine_rom(616);
     when "001001101001" => data <= sine_rom(617);
     when "001001101010" => data <= sine_rom(618);
     when "001001101011" => data <= sine_rom(619);
     when "001001101100" => data <= sine_rom(620);
     when "001001101101" => data <= sine_rom(621);
     when "001001101110" => data <= sine_rom(622);
     when "001001101111" => data <= sine_rom(623);
     when "001001110000" => data <= sine_rom(624);
     when "001001110001" => data <= sine_rom(625);
     when "001001110010" => data <= sine_rom(626);
     when "001001110011" => data <= sine_rom(627);
     when "001001110100" => data <= sine_rom(628);
     when "001001110101" => data <= sine_rom(629);
     when "001001110110" => data <= sine_rom(630);
     when "001001110111" => data <= sine_rom(631);
     when "001001111000" => data <= sine_rom(632);
     when "001001111001" => data <= sine_rom(633);
     when "001001111010" => data <= sine_rom(634);
     when "001001111011" => data <= sine_rom(635);
     when "001001111100" => data <= sine_rom(636);
     when "001001111101" => data <= sine_rom(637);
     when "001001111110" => data <= sine_rom(638);
     when "001001111111" => data <= sine_rom(639);
     when "001010000000" => data <= sine_rom(640);
     when "001010000001" => data <= sine_rom(641);
     when "001010000010" => data <= sine_rom(642);
     when "001010000011" => data <= sine_rom(643);
     when "001010000100" => data <= sine_rom(644);
     when "001010000101" => data <= sine_rom(645);
     when "001010000110" => data <= sine_rom(646);
     when "001010000111" => data <= sine_rom(647);
     when "001010001000" => data <= sine_rom(648);
     when "001010001001" => data <= sine_rom(649);
     when "001010001010" => data <= sine_rom(650);
     when "001010001011" => data <= sine_rom(651);
     when "001010001100" => data <= sine_rom(652);
     when "001010001101" => data <= sine_rom(653);
     when "001010001110" => data <= sine_rom(654);
     when "001010001111" => data <= sine_rom(655);
     when "001010010000" => data <= sine_rom(656);
     when "001010010001" => data <= sine_rom(657);
     when "001010010010" => data <= sine_rom(658);
     when "001010010011" => data <= sine_rom(659);
     when "001010010100" => data <= sine_rom(660);
     when "001010010101" => data <= sine_rom(661);
     when "001010010110" => data <= sine_rom(662);
     when "001010010111" => data <= sine_rom(663);
     when "001010011000" => data <= sine_rom(664);
     when "001010011001" => data <= sine_rom(665);
     when "001010011010" => data <= sine_rom(666);
     when "001010011011" => data <= sine_rom(667);
     when "001010011100" => data <= sine_rom(668);
     when "001010011101" => data <= sine_rom(669);
     when "001010011110" => data <= sine_rom(670);
     when "001010011111" => data <= sine_rom(671);
     when "001010100000" => data <= sine_rom(672);
     when "001010100001" => data <= sine_rom(673);
     when "001010100010" => data <= sine_rom(674);
     when "001010100011" => data <= sine_rom(675);
     when "001010100100" => data <= sine_rom(676);
     when "001010100101" => data <= sine_rom(677);
     when "001010100110" => data <= sine_rom(678);
     when "001010100111" => data <= sine_rom(679);
     when "001010101000" => data <= sine_rom(680);
     when "001010101001" => data <= sine_rom(681);
     when "001010101010" => data <= sine_rom(682);
     when "001010101011" => data <= sine_rom(683);
     when "001010101100" => data <= sine_rom(684);
     when "001010101101" => data <= sine_rom(685);
     when "001010101110" => data <= sine_rom(686);
     when "001010101111" => data <= sine_rom(687);
     when "001010110000" => data <= sine_rom(688);
     when "001010110001" => data <= sine_rom(689);
     when "001010110010" => data <= sine_rom(690);
     when "001010110011" => data <= sine_rom(691);
     when "001010110100" => data <= sine_rom(692);
     when "001010110101" => data <= sine_rom(693);
     when "001010110110" => data <= sine_rom(694);
     when "001010110111" => data <= sine_rom(695);
     when "001010111000" => data <= sine_rom(696);
     when "001010111001" => data <= sine_rom(697);
     when "001010111010" => data <= sine_rom(698);
     when "001010111011" => data <= sine_rom(699);
     when "001010111100" => data <= sine_rom(700);
     when "001010111101" => data <= sine_rom(701);
     when "001010111110" => data <= sine_rom(702);
     when "001010111111" => data <= sine_rom(703);
     when "001011000000" => data <= sine_rom(704);
     when "001011000001" => data <= sine_rom(705);
     when "001011000010" => data <= sine_rom(706);
     when "001011000011" => data <= sine_rom(707);
     when "001011000100" => data <= sine_rom(708);
     when "001011000101" => data <= sine_rom(709);
     when "001011000110" => data <= sine_rom(710);
     when "001011000111" => data <= sine_rom(711);
     when "001011001000" => data <= sine_rom(712);
     when "001011001001" => data <= sine_rom(713);
     when "001011001010" => data <= sine_rom(714);
     when "001011001011" => data <= sine_rom(715);
     when "001011001100" => data <= sine_rom(716);
     when "001011001101" => data <= sine_rom(717);
     when "001011001110" => data <= sine_rom(718);
     when "001011001111" => data <= sine_rom(719);
     when "001011010000" => data <= sine_rom(720);
     when "001011010001" => data <= sine_rom(721);
     when "001011010010" => data <= sine_rom(722);
     when "001011010011" => data <= sine_rom(723);
     when "001011010100" => data <= sine_rom(724);
     when "001011010101" => data <= sine_rom(725);
     when "001011010110" => data <= sine_rom(726);
     when "001011010111" => data <= sine_rom(727);
     when "001011011000" => data <= sine_rom(728);
     when "001011011001" => data <= sine_rom(729);
     when "001011011010" => data <= sine_rom(730);
     when "001011011011" => data <= sine_rom(731);
     when "001011011100" => data <= sine_rom(732);
     when "001011011101" => data <= sine_rom(733);
     when "001011011110" => data <= sine_rom(734);
     when "001011011111" => data <= sine_rom(735);
     when "001011100000" => data <= sine_rom(736);
     when "001011100001" => data <= sine_rom(737);
     when "001011100010" => data <= sine_rom(738);
     when "001011100011" => data <= sine_rom(739);
     when "001011100100" => data <= sine_rom(740);
     when "001011100101" => data <= sine_rom(741);
     when "001011100110" => data <= sine_rom(742);
     when "001011100111" => data <= sine_rom(743);
     when "001011101000" => data <= sine_rom(744);
     when "001011101001" => data <= sine_rom(745);
     when "001011101010" => data <= sine_rom(746);
     when "001011101011" => data <= sine_rom(747);
     when "001011101100" => data <= sine_rom(748);
     when "001011101101" => data <= sine_rom(749);
     when "001011101110" => data <= sine_rom(750);
     when "001011101111" => data <= sine_rom(751);
     when "001011110000" => data <= sine_rom(752);
     when "001011110001" => data <= sine_rom(753);
     when "001011110010" => data <= sine_rom(754);
     when "001011110011" => data <= sine_rom(755);
     when "001011110100" => data <= sine_rom(756);
     when "001011110101" => data <= sine_rom(757);
     when "001011110110" => data <= sine_rom(758);
     when "001011110111" => data <= sine_rom(759);
     when "001011111000" => data <= sine_rom(760);
     when "001011111001" => data <= sine_rom(761);
     when "001011111010" => data <= sine_rom(762);
     when "001011111011" => data <= sine_rom(763);
     when "001011111100" => data <= sine_rom(764);
     when "001011111101" => data <= sine_rom(765);
     when "001011111110" => data <= sine_rom(766);
     when "001011111111" => data <= sine_rom(767);
     when "001100000000" => data <= sine_rom(768);
     when "001100000001" => data <= sine_rom(769);
     when "001100000010" => data <= sine_rom(770);
     when "001100000011" => data <= sine_rom(771);
     when "001100000100" => data <= sine_rom(772);
     when "001100000101" => data <= sine_rom(773);
     when "001100000110" => data <= sine_rom(774);
     when "001100000111" => data <= sine_rom(775);
     when "001100001000" => data <= sine_rom(776);
     when "001100001001" => data <= sine_rom(777);
     when "001100001010" => data <= sine_rom(778);
     when "001100001011" => data <= sine_rom(779);
     when "001100001100" => data <= sine_rom(780);
     when "001100001101" => data <= sine_rom(781);
     when "001100001110" => data <= sine_rom(782);
     when "001100001111" => data <= sine_rom(783);
     when "001100010000" => data <= sine_rom(784);
     when "001100010001" => data <= sine_rom(785);
     when "001100010010" => data <= sine_rom(786);
     when "001100010011" => data <= sine_rom(787);
     when "001100010100" => data <= sine_rom(788);
     when "001100010101" => data <= sine_rom(789);
     when "001100010110" => data <= sine_rom(790);
     when "001100010111" => data <= sine_rom(791);
     when "001100011000" => data <= sine_rom(792);
     when "001100011001" => data <= sine_rom(793);
     when "001100011010" => data <= sine_rom(794);
     when "001100011011" => data <= sine_rom(795);
     when "001100011100" => data <= sine_rom(796);
     when "001100011101" => data <= sine_rom(797);
     when "001100011110" => data <= sine_rom(798);
     when "001100011111" => data <= sine_rom(799);
     when "001100100000" => data <= sine_rom(800);
     when "001100100001" => data <= sine_rom(801);
     when "001100100010" => data <= sine_rom(802);
     when "001100100011" => data <= sine_rom(803);
     when "001100100100" => data <= sine_rom(804);
     when "001100100101" => data <= sine_rom(805);
     when "001100100110" => data <= sine_rom(806);
     when "001100100111" => data <= sine_rom(807);
     when "001100101000" => data <= sine_rom(808);
     when "001100101001" => data <= sine_rom(809);
     when "001100101010" => data <= sine_rom(810);
     when "001100101011" => data <= sine_rom(811);
     when "001100101100" => data <= sine_rom(812);
     when "001100101101" => data <= sine_rom(813);
     when "001100101110" => data <= sine_rom(814);
     when "001100101111" => data <= sine_rom(815);
     when "001100110000" => data <= sine_rom(816);
     when "001100110001" => data <= sine_rom(817);
     when "001100110010" => data <= sine_rom(818);
     when "001100110011" => data <= sine_rom(819);
     when "001100110100" => data <= sine_rom(820);
     when "001100110101" => data <= sine_rom(821);
     when "001100110110" => data <= sine_rom(822);
     when "001100110111" => data <= sine_rom(823);
     when "001100111000" => data <= sine_rom(824);
     when "001100111001" => data <= sine_rom(825);
     when "001100111010" => data <= sine_rom(826);
     when "001100111011" => data <= sine_rom(827);
     when "001100111100" => data <= sine_rom(828);
     when "001100111101" => data <= sine_rom(829);
     when "001100111110" => data <= sine_rom(830);
     when "001100111111" => data <= sine_rom(831);
     when "001101000000" => data <= sine_rom(832);
     when "001101000001" => data <= sine_rom(833);
     when "001101000010" => data <= sine_rom(834);
     when "001101000011" => data <= sine_rom(835);
     when "001101000100" => data <= sine_rom(836);
     when "001101000101" => data <= sine_rom(837);
     when "001101000110" => data <= sine_rom(838);
     when "001101000111" => data <= sine_rom(839);
     when "001101001000" => data <= sine_rom(840);
     when "001101001001" => data <= sine_rom(841);
     when "001101001010" => data <= sine_rom(842);
     when "001101001011" => data <= sine_rom(843);
     when "001101001100" => data <= sine_rom(844);
     when "001101001101" => data <= sine_rom(845);
     when "001101001110" => data <= sine_rom(846);
     when "001101001111" => data <= sine_rom(847);
     when "001101010000" => data <= sine_rom(848);
     when "001101010001" => data <= sine_rom(849);
     when "001101010010" => data <= sine_rom(850);
     when "001101010011" => data <= sine_rom(851);
     when "001101010100" => data <= sine_rom(852);
     when "001101010101" => data <= sine_rom(853);
     when "001101010110" => data <= sine_rom(854);
     when "001101010111" => data <= sine_rom(855);
     when "001101011000" => data <= sine_rom(856);
     when "001101011001" => data <= sine_rom(857);
     when "001101011010" => data <= sine_rom(858);
     when "001101011011" => data <= sine_rom(859);
     when "001101011100" => data <= sine_rom(860);
     when "001101011101" => data <= sine_rom(861);
     when "001101011110" => data <= sine_rom(862);
     when "001101011111" => data <= sine_rom(863);
     when "001101100000" => data <= sine_rom(864);
     when "001101100001" => data <= sine_rom(865);
     when "001101100010" => data <= sine_rom(866);
     when "001101100011" => data <= sine_rom(867);
     when "001101100100" => data <= sine_rom(868);
     when "001101100101" => data <= sine_rom(869);
     when "001101100110" => data <= sine_rom(870);
     when "001101100111" => data <= sine_rom(871);
     when "001101101000" => data <= sine_rom(872);
     when "001101101001" => data <= sine_rom(873);
     when "001101101010" => data <= sine_rom(874);
     when "001101101011" => data <= sine_rom(875);
     when "001101101100" => data <= sine_rom(876);
     when "001101101101" => data <= sine_rom(877);
     when "001101101110" => data <= sine_rom(878);
     when "001101101111" => data <= sine_rom(879);
     when "001101110000" => data <= sine_rom(880);
     when "001101110001" => data <= sine_rom(881);
     when "001101110010" => data <= sine_rom(882);
     when "001101110011" => data <= sine_rom(883);
     when "001101110100" => data <= sine_rom(884);
     when "001101110101" => data <= sine_rom(885);
     when "001101110110" => data <= sine_rom(886);
     when "001101110111" => data <= sine_rom(887);
     when "001101111000" => data <= sine_rom(888);
     when "001101111001" => data <= sine_rom(889);
     when "001101111010" => data <= sine_rom(890);
     when "001101111011" => data <= sine_rom(891);
     when "001101111100" => data <= sine_rom(892);
     when "001101111101" => data <= sine_rom(893);
     when "001101111110" => data <= sine_rom(894);
     when "001101111111" => data <= sine_rom(895);
     when "001110000000" => data <= sine_rom(896);
     when "001110000001" => data <= sine_rom(897);
     when "001110000010" => data <= sine_rom(898);
     when "001110000011" => data <= sine_rom(899);
     when "001110000100" => data <= sine_rom(900);
     when "001110000101" => data <= sine_rom(901);
     when "001110000110" => data <= sine_rom(902);
     when "001110000111" => data <= sine_rom(903);
     when "001110001000" => data <= sine_rom(904);
     when "001110001001" => data <= sine_rom(905);
     when "001110001010" => data <= sine_rom(906);
     when "001110001011" => data <= sine_rom(907);
     when "001110001100" => data <= sine_rom(908);
     when "001110001101" => data <= sine_rom(909);
     when "001110001110" => data <= sine_rom(910);
     when "001110001111" => data <= sine_rom(911);
     when "001110010000" => data <= sine_rom(912);
     when "001110010001" => data <= sine_rom(913);
     when "001110010010" => data <= sine_rom(914);
     when "001110010011" => data <= sine_rom(915);
     when "001110010100" => data <= sine_rom(916);
     when "001110010101" => data <= sine_rom(917);
     when "001110010110" => data <= sine_rom(918);
     when "001110010111" => data <= sine_rom(919);
     when "001110011000" => data <= sine_rom(920);
     when "001110011001" => data <= sine_rom(921);
     when "001110011010" => data <= sine_rom(922);
     when "001110011011" => data <= sine_rom(923);
     when "001110011100" => data <= sine_rom(924);
     when "001110011101" => data <= sine_rom(925);
     when "001110011110" => data <= sine_rom(926);
     when "001110011111" => data <= sine_rom(927);
     when "001110100000" => data <= sine_rom(928);
     when "001110100001" => data <= sine_rom(929);
     when "001110100010" => data <= sine_rom(930);
     when "001110100011" => data <= sine_rom(931);
     when "001110100100" => data <= sine_rom(932);
     when "001110100101" => data <= sine_rom(933);
     when "001110100110" => data <= sine_rom(934);
     when "001110100111" => data <= sine_rom(935);
     when "001110101000" => data <= sine_rom(936);
     when "001110101001" => data <= sine_rom(937);
     when "001110101010" => data <= sine_rom(938);
     when "001110101011" => data <= sine_rom(939);
     when "001110101100" => data <= sine_rom(940);
     when "001110101101" => data <= sine_rom(941);
     when "001110101110" => data <= sine_rom(942);
     when "001110101111" => data <= sine_rom(943);
     when "001110110000" => data <= sine_rom(944);
     when "001110110001" => data <= sine_rom(945);
     when "001110110010" => data <= sine_rom(946);
     when "001110110011" => data <= sine_rom(947);
     when "001110110100" => data <= sine_rom(948);
     when "001110110101" => data <= sine_rom(949);
     when "001110110110" => data <= sine_rom(950);
     when "001110110111" => data <= sine_rom(951);
     when "001110111000" => data <= sine_rom(952);
     when "001110111001" => data <= sine_rom(953);
     when "001110111010" => data <= sine_rom(954);
     when "001110111011" => data <= sine_rom(955);
     when "001110111100" => data <= sine_rom(956);
     when "001110111101" => data <= sine_rom(957);
     when "001110111110" => data <= sine_rom(958);
     when "001110111111" => data <= sine_rom(959);
     when "001111000000" => data <= sine_rom(960);
     when "001111000001" => data <= sine_rom(961);
     when "001111000010" => data <= sine_rom(962);
     when "001111000011" => data <= sine_rom(963);
     when "001111000100" => data <= sine_rom(964);
     when "001111000101" => data <= sine_rom(965);
     when "001111000110" => data <= sine_rom(966);
     when "001111000111" => data <= sine_rom(967);
     when "001111001000" => data <= sine_rom(968);
     when "001111001001" => data <= sine_rom(969);
     when "001111001010" => data <= sine_rom(970);
     when "001111001011" => data <= sine_rom(971);
     when "001111001100" => data <= sine_rom(972);
     when "001111001101" => data <= sine_rom(973);
     when "001111001110" => data <= sine_rom(974);
     when "001111001111" => data <= sine_rom(975);
     when "001111010000" => data <= sine_rom(976);
     when "001111010001" => data <= sine_rom(977);
     when "001111010010" => data <= sine_rom(978);
     when "001111010011" => data <= sine_rom(979);
     when "001111010100" => data <= sine_rom(980);
     when "001111010101" => data <= sine_rom(981);
     when "001111010110" => data <= sine_rom(982);
     when "001111010111" => data <= sine_rom(983);
     when "001111011000" => data <= sine_rom(984);
     when "001111011001" => data <= sine_rom(985);
     when "001111011010" => data <= sine_rom(986);
     when "001111011011" => data <= sine_rom(987);
     when "001111011100" => data <= sine_rom(988);
     when "001111011101" => data <= sine_rom(989);
     when "001111011110" => data <= sine_rom(990);
     when "001111011111" => data <= sine_rom(991);
     when "001111100000" => data <= sine_rom(992);
     when "001111100001" => data <= sine_rom(993);
     when "001111100010" => data <= sine_rom(994);
     when "001111100011" => data <= sine_rom(995);
     when "001111100100" => data <= sine_rom(996);
     when "001111100101" => data <= sine_rom(997);
     when "001111100110" => data <= sine_rom(998);
     when "001111100111" => data <= sine_rom(999);
     when "001111101000" => data <= sine_rom(1000);
     when "001111101001" => data <= sine_rom(1001);
     when "001111101010" => data <= sine_rom(1002);
     when "001111101011" => data <= sine_rom(1003);
     when "001111101100" => data <= sine_rom(1004);
     when "001111101101" => data <= sine_rom(1005);
     when "001111101110" => data <= sine_rom(1006);
     when "001111101111" => data <= sine_rom(1007);
     when "001111110000" => data <= sine_rom(1008);
     when "001111110001" => data <= sine_rom(1009);
     when "001111110010" => data <= sine_rom(1010);
     when "001111110011" => data <= sine_rom(1011);
     when "001111110100" => data <= sine_rom(1012);
     when "001111110101" => data <= sine_rom(1013);
     when "001111110110" => data <= sine_rom(1014);
     when "001111110111" => data <= sine_rom(1015);
     when "001111111000" => data <= sine_rom(1016);
     when "001111111001" => data <= sine_rom(1017);
     when "001111111010" => data <= sine_rom(1018);
     when "001111111011" => data <= sine_rom(1019);
     when "001111111100" => data <= sine_rom(1020);
     when "001111111101" => data <= sine_rom(1021);
     when "001111111110" => data <= sine_rom(1022);
     when "001111111111" => data <= sine_rom(1023);
     when "010000000000" => data <= sine_rom(1024);
     when "010000000001" => data <= sine_rom(1025);
     when "010000000010" => data <= sine_rom(1026);
     when "010000000011" => data <= sine_rom(1027);
     when "010000000100" => data <= sine_rom(1028);
     when "010000000101" => data <= sine_rom(1029);
     when "010000000110" => data <= sine_rom(1030);
     when "010000000111" => data <= sine_rom(1031);
     when "010000001000" => data <= sine_rom(1032);
     when "010000001001" => data <= sine_rom(1033);
     when "010000001010" => data <= sine_rom(1034);
     when "010000001011" => data <= sine_rom(1035);
     when "010000001100" => data <= sine_rom(1036);
     when "010000001101" => data <= sine_rom(1037);
     when "010000001110" => data <= sine_rom(1038);
     when "010000001111" => data <= sine_rom(1039);
     when "010000010000" => data <= sine_rom(1040);
     when "010000010001" => data <= sine_rom(1041);
     when "010000010010" => data <= sine_rom(1042);
     when "010000010011" => data <= sine_rom(1043);
     when "010000010100" => data <= sine_rom(1044);
     when "010000010101" => data <= sine_rom(1045);
     when "010000010110" => data <= sine_rom(1046);
     when "010000010111" => data <= sine_rom(1047);
     when "010000011000" => data <= sine_rom(1048);
     when "010000011001" => data <= sine_rom(1049);
     when "010000011010" => data <= sine_rom(1050);
     when "010000011011" => data <= sine_rom(1051);
     when "010000011100" => data <= sine_rom(1052);
     when "010000011101" => data <= sine_rom(1053);
     when "010000011110" => data <= sine_rom(1054);
     when "010000011111" => data <= sine_rom(1055);
     when "010000100000" => data <= sine_rom(1056);
     when "010000100001" => data <= sine_rom(1057);
     when "010000100010" => data <= sine_rom(1058);
     when "010000100011" => data <= sine_rom(1059);
     when "010000100100" => data <= sine_rom(1060);
     when "010000100101" => data <= sine_rom(1061);
     when "010000100110" => data <= sine_rom(1062);
     when "010000100111" => data <= sine_rom(1063);
     when "010000101000" => data <= sine_rom(1064);
     when "010000101001" => data <= sine_rom(1065);
     when "010000101010" => data <= sine_rom(1066);
     when "010000101011" => data <= sine_rom(1067);
     when "010000101100" => data <= sine_rom(1068);
     when "010000101101" => data <= sine_rom(1069);
     when "010000101110" => data <= sine_rom(1070);
     when "010000101111" => data <= sine_rom(1071);
     when "010000110000" => data <= sine_rom(1072);
     when "010000110001" => data <= sine_rom(1073);
     when "010000110010" => data <= sine_rom(1074);
     when "010000110011" => data <= sine_rom(1075);
     when "010000110100" => data <= sine_rom(1076);
     when "010000110101" => data <= sine_rom(1077);
     when "010000110110" => data <= sine_rom(1078);
     when "010000110111" => data <= sine_rom(1079);
     when "010000111000" => data <= sine_rom(1080);
     when "010000111001" => data <= sine_rom(1081);
     when "010000111010" => data <= sine_rom(1082);
     when "010000111011" => data <= sine_rom(1083);
     when "010000111100" => data <= sine_rom(1084);
     when "010000111101" => data <= sine_rom(1085);
     when "010000111110" => data <= sine_rom(1086);
     when "010000111111" => data <= sine_rom(1087);
     when "010001000000" => data <= sine_rom(1088);
     when "010001000001" => data <= sine_rom(1089);
     when "010001000010" => data <= sine_rom(1090);
     when "010001000011" => data <= sine_rom(1091);
     when "010001000100" => data <= sine_rom(1092);
     when "010001000101" => data <= sine_rom(1093);
     when "010001000110" => data <= sine_rom(1094);
     when "010001000111" => data <= sine_rom(1095);
     when "010001001000" => data <= sine_rom(1096);
     when "010001001001" => data <= sine_rom(1097);
     when "010001001010" => data <= sine_rom(1098);
     when "010001001011" => data <= sine_rom(1099);
     when "010001001100" => data <= sine_rom(1100);
     when "010001001101" => data <= sine_rom(1101);
     when "010001001110" => data <= sine_rom(1102);
     when "010001001111" => data <= sine_rom(1103);
     when "010001010000" => data <= sine_rom(1104);
     when "010001010001" => data <= sine_rom(1105);
     when "010001010010" => data <= sine_rom(1106);
     when "010001010011" => data <= sine_rom(1107);
     when "010001010100" => data <= sine_rom(1108);
     when "010001010101" => data <= sine_rom(1109);
     when "010001010110" => data <= sine_rom(1110);
     when "010001010111" => data <= sine_rom(1111);
     when "010001011000" => data <= sine_rom(1112);
     when "010001011001" => data <= sine_rom(1113);
     when "010001011010" => data <= sine_rom(1114);
     when "010001011011" => data <= sine_rom(1115);
     when "010001011100" => data <= sine_rom(1116);
     when "010001011101" => data <= sine_rom(1117);
     when "010001011110" => data <= sine_rom(1118);
     when "010001011111" => data <= sine_rom(1119);
     when "010001100000" => data <= sine_rom(1120);
     when "010001100001" => data <= sine_rom(1121);
     when "010001100010" => data <= sine_rom(1122);
     when "010001100011" => data <= sine_rom(1123);
     when "010001100100" => data <= sine_rom(1124);
     when "010001100101" => data <= sine_rom(1125);
     when "010001100110" => data <= sine_rom(1126);
     when "010001100111" => data <= sine_rom(1127);
     when "010001101000" => data <= sine_rom(1128);
     when "010001101001" => data <= sine_rom(1129);
     when "010001101010" => data <= sine_rom(1130);
     when "010001101011" => data <= sine_rom(1131);
     when "010001101100" => data <= sine_rom(1132);
     when "010001101101" => data <= sine_rom(1133);
     when "010001101110" => data <= sine_rom(1134);
     when "010001101111" => data <= sine_rom(1135);
     when "010001110000" => data <= sine_rom(1136);
     when "010001110001" => data <= sine_rom(1137);
     when "010001110010" => data <= sine_rom(1138);
     when "010001110011" => data <= sine_rom(1139);
     when "010001110100" => data <= sine_rom(1140);
     when "010001110101" => data <= sine_rom(1141);
     when "010001110110" => data <= sine_rom(1142);
     when "010001110111" => data <= sine_rom(1143);
     when "010001111000" => data <= sine_rom(1144);
     when "010001111001" => data <= sine_rom(1145);
     when "010001111010" => data <= sine_rom(1146);
     when "010001111011" => data <= sine_rom(1147);
     when "010001111100" => data <= sine_rom(1148);
     when "010001111101" => data <= sine_rom(1149);
     when "010001111110" => data <= sine_rom(1150);
     when "010001111111" => data <= sine_rom(1151);
     when "010010000000" => data <= sine_rom(1152);
     when "010010000001" => data <= sine_rom(1153);
     when "010010000010" => data <= sine_rom(1154);
     when "010010000011" => data <= sine_rom(1155);
     when "010010000100" => data <= sine_rom(1156);
     when "010010000101" => data <= sine_rom(1157);
     when "010010000110" => data <= sine_rom(1158);
     when "010010000111" => data <= sine_rom(1159);
     when "010010001000" => data <= sine_rom(1160);
     when "010010001001" => data <= sine_rom(1161);
     when "010010001010" => data <= sine_rom(1162);
     when "010010001011" => data <= sine_rom(1163);
     when "010010001100" => data <= sine_rom(1164);
     when "010010001101" => data <= sine_rom(1165);
     when "010010001110" => data <= sine_rom(1166);
     when "010010001111" => data <= sine_rom(1167);
     when "010010010000" => data <= sine_rom(1168);
     when "010010010001" => data <= sine_rom(1169);
     when "010010010010" => data <= sine_rom(1170);
     when "010010010011" => data <= sine_rom(1171);
     when "010010010100" => data <= sine_rom(1172);
     when "010010010101" => data <= sine_rom(1173);
     when "010010010110" => data <= sine_rom(1174);
     when "010010010111" => data <= sine_rom(1175);
     when "010010011000" => data <= sine_rom(1176);
     when "010010011001" => data <= sine_rom(1177);
     when "010010011010" => data <= sine_rom(1178);
     when "010010011011" => data <= sine_rom(1179);
     when "010010011100" => data <= sine_rom(1180);
     when "010010011101" => data <= sine_rom(1181);
     when "010010011110" => data <= sine_rom(1182);
     when "010010011111" => data <= sine_rom(1183);
     when "010010100000" => data <= sine_rom(1184);
     when "010010100001" => data <= sine_rom(1185);
     when "010010100010" => data <= sine_rom(1186);
     when "010010100011" => data <= sine_rom(1187);
     when "010010100100" => data <= sine_rom(1188);
     when "010010100101" => data <= sine_rom(1189);
     when "010010100110" => data <= sine_rom(1190);
     when "010010100111" => data <= sine_rom(1191);
     when "010010101000" => data <= sine_rom(1192);
     when "010010101001" => data <= sine_rom(1193);
     when "010010101010" => data <= sine_rom(1194);
     when "010010101011" => data <= sine_rom(1195);
     when "010010101100" => data <= sine_rom(1196);
     when "010010101101" => data <= sine_rom(1197);
     when "010010101110" => data <= sine_rom(1198);
     when "010010101111" => data <= sine_rom(1199);
     when "010010110000" => data <= sine_rom(1200);
     when "010010110001" => data <= sine_rom(1201);
     when "010010110010" => data <= sine_rom(1202);
     when "010010110011" => data <= sine_rom(1203);
     when "010010110100" => data <= sine_rom(1204);
     when "010010110101" => data <= sine_rom(1205);
     when "010010110110" => data <= sine_rom(1206);
     when "010010110111" => data <= sine_rom(1207);
     when "010010111000" => data <= sine_rom(1208);
     when "010010111001" => data <= sine_rom(1209);
     when "010010111010" => data <= sine_rom(1210);
     when "010010111011" => data <= sine_rom(1211);
     when "010010111100" => data <= sine_rom(1212);
     when "010010111101" => data <= sine_rom(1213);
     when "010010111110" => data <= sine_rom(1214);
     when "010010111111" => data <= sine_rom(1215);
     when "010011000000" => data <= sine_rom(1216);
     when "010011000001" => data <= sine_rom(1217);
     when "010011000010" => data <= sine_rom(1218);
     when "010011000011" => data <= sine_rom(1219);
     when "010011000100" => data <= sine_rom(1220);
     when "010011000101" => data <= sine_rom(1221);
     when "010011000110" => data <= sine_rom(1222);
     when "010011000111" => data <= sine_rom(1223);
     when "010011001000" => data <= sine_rom(1224);
     when "010011001001" => data <= sine_rom(1225);
     when "010011001010" => data <= sine_rom(1226);
     when "010011001011" => data <= sine_rom(1227);
     when "010011001100" => data <= sine_rom(1228);
     when "010011001101" => data <= sine_rom(1229);
     when "010011001110" => data <= sine_rom(1230);
     when "010011001111" => data <= sine_rom(1231);
     when "010011010000" => data <= sine_rom(1232);
     when "010011010001" => data <= sine_rom(1233);
     when "010011010010" => data <= sine_rom(1234);
     when "010011010011" => data <= sine_rom(1235);
     when "010011010100" => data <= sine_rom(1236);
     when "010011010101" => data <= sine_rom(1237);
     when "010011010110" => data <= sine_rom(1238);
     when "010011010111" => data <= sine_rom(1239);
     when "010011011000" => data <= sine_rom(1240);
     when "010011011001" => data <= sine_rom(1241);
     when "010011011010" => data <= sine_rom(1242);
     when "010011011011" => data <= sine_rom(1243);
     when "010011011100" => data <= sine_rom(1244);
     when "010011011101" => data <= sine_rom(1245);
     when "010011011110" => data <= sine_rom(1246);
     when "010011011111" => data <= sine_rom(1247);
     when "010011100000" => data <= sine_rom(1248);
     when "010011100001" => data <= sine_rom(1249);
     when "010011100010" => data <= sine_rom(1250);
     when "010011100011" => data <= sine_rom(1251);
     when "010011100100" => data <= sine_rom(1252);
     when "010011100101" => data <= sine_rom(1253);
     when "010011100110" => data <= sine_rom(1254);
     when "010011100111" => data <= sine_rom(1255);
     when "010011101000" => data <= sine_rom(1256);
     when "010011101001" => data <= sine_rom(1257);
     when "010011101010" => data <= sine_rom(1258);
     when "010011101011" => data <= sine_rom(1259);
     when "010011101100" => data <= sine_rom(1260);
     when "010011101101" => data <= sine_rom(1261);
     when "010011101110" => data <= sine_rom(1262);
     when "010011101111" => data <= sine_rom(1263);
     when "010011110000" => data <= sine_rom(1264);
     when "010011110001" => data <= sine_rom(1265);
     when "010011110010" => data <= sine_rom(1266);
     when "010011110011" => data <= sine_rom(1267);
     when "010011110100" => data <= sine_rom(1268);
     when "010011110101" => data <= sine_rom(1269);
     when "010011110110" => data <= sine_rom(1270);
     when "010011110111" => data <= sine_rom(1271);
     when "010011111000" => data <= sine_rom(1272);
     when "010011111001" => data <= sine_rom(1273);
     when "010011111010" => data <= sine_rom(1274);
     when "010011111011" => data <= sine_rom(1275);
     when "010011111100" => data <= sine_rom(1276);
     when "010011111101" => data <= sine_rom(1277);
     when "010011111110" => data <= sine_rom(1278);
     when "010011111111" => data <= sine_rom(1279);
     when "010100000000" => data <= sine_rom(1280);
     when "010100000001" => data <= sine_rom(1281);
     when "010100000010" => data <= sine_rom(1282);
     when "010100000011" => data <= sine_rom(1283);
     when "010100000100" => data <= sine_rom(1284);
     when "010100000101" => data <= sine_rom(1285);
     when "010100000110" => data <= sine_rom(1286);
     when "010100000111" => data <= sine_rom(1287);
     when "010100001000" => data <= sine_rom(1288);
     when "010100001001" => data <= sine_rom(1289);
     when "010100001010" => data <= sine_rom(1290);
     when "010100001011" => data <= sine_rom(1291);
     when "010100001100" => data <= sine_rom(1292);
     when "010100001101" => data <= sine_rom(1293);
     when "010100001110" => data <= sine_rom(1294);
     when "010100001111" => data <= sine_rom(1295);
     when "010100010000" => data <= sine_rom(1296);
     when "010100010001" => data <= sine_rom(1297);
     when "010100010010" => data <= sine_rom(1298);
     when "010100010011" => data <= sine_rom(1299);
     when "010100010100" => data <= sine_rom(1300);
     when "010100010101" => data <= sine_rom(1301);
     when "010100010110" => data <= sine_rom(1302);
     when "010100010111" => data <= sine_rom(1303);
     when "010100011000" => data <= sine_rom(1304);
     when "010100011001" => data <= sine_rom(1305);
     when "010100011010" => data <= sine_rom(1306);
     when "010100011011" => data <= sine_rom(1307);
     when "010100011100" => data <= sine_rom(1308);
     when "010100011101" => data <= sine_rom(1309);
     when "010100011110" => data <= sine_rom(1310);
     when "010100011111" => data <= sine_rom(1311);
     when "010100100000" => data <= sine_rom(1312);
     when "010100100001" => data <= sine_rom(1313);
     when "010100100010" => data <= sine_rom(1314);
     when "010100100011" => data <= sine_rom(1315);
     when "010100100100" => data <= sine_rom(1316);
     when "010100100101" => data <= sine_rom(1317);
     when "010100100110" => data <= sine_rom(1318);
     when "010100100111" => data <= sine_rom(1319);
     when "010100101000" => data <= sine_rom(1320);
     when "010100101001" => data <= sine_rom(1321);
     when "010100101010" => data <= sine_rom(1322);
     when "010100101011" => data <= sine_rom(1323);
     when "010100101100" => data <= sine_rom(1324);
     when "010100101101" => data <= sine_rom(1325);
     when "010100101110" => data <= sine_rom(1326);
     when "010100101111" => data <= sine_rom(1327);
     when "010100110000" => data <= sine_rom(1328);
     when "010100110001" => data <= sine_rom(1329);
     when "010100110010" => data <= sine_rom(1330);
     when "010100110011" => data <= sine_rom(1331);
     when "010100110100" => data <= sine_rom(1332);
     when "010100110101" => data <= sine_rom(1333);
     when "010100110110" => data <= sine_rom(1334);
     when "010100110111" => data <= sine_rom(1335);
     when "010100111000" => data <= sine_rom(1336);
     when "010100111001" => data <= sine_rom(1337);
     when "010100111010" => data <= sine_rom(1338);
     when "010100111011" => data <= sine_rom(1339);
     when "010100111100" => data <= sine_rom(1340);
     when "010100111101" => data <= sine_rom(1341);
     when "010100111110" => data <= sine_rom(1342);
     when "010100111111" => data <= sine_rom(1343);
     when "010101000000" => data <= sine_rom(1344);
     when "010101000001" => data <= sine_rom(1345);
     when "010101000010" => data <= sine_rom(1346);
     when "010101000011" => data <= sine_rom(1347);
     when "010101000100" => data <= sine_rom(1348);
     when "010101000101" => data <= sine_rom(1349);
     when "010101000110" => data <= sine_rom(1350);
     when "010101000111" => data <= sine_rom(1351);
     when "010101001000" => data <= sine_rom(1352);
     when "010101001001" => data <= sine_rom(1353);
     when "010101001010" => data <= sine_rom(1354);
     when "010101001011" => data <= sine_rom(1355);
     when "010101001100" => data <= sine_rom(1356);
     when "010101001101" => data <= sine_rom(1357);
     when "010101001110" => data <= sine_rom(1358);
     when "010101001111" => data <= sine_rom(1359);
     when "010101010000" => data <= sine_rom(1360);
     when "010101010001" => data <= sine_rom(1361);
     when "010101010010" => data <= sine_rom(1362);
     when "010101010011" => data <= sine_rom(1363);
     when "010101010100" => data <= sine_rom(1364);
     when "010101010101" => data <= sine_rom(1365);
     when "010101010110" => data <= sine_rom(1366);
     when "010101010111" => data <= sine_rom(1367);
     when "010101011000" => data <= sine_rom(1368);
     when "010101011001" => data <= sine_rom(1369);
     when "010101011010" => data <= sine_rom(1370);
     when "010101011011" => data <= sine_rom(1371);
     when "010101011100" => data <= sine_rom(1372);
     when "010101011101" => data <= sine_rom(1373);
     when "010101011110" => data <= sine_rom(1374);
     when "010101011111" => data <= sine_rom(1375);
     when "010101100000" => data <= sine_rom(1376);
     when "010101100001" => data <= sine_rom(1377);
     when "010101100010" => data <= sine_rom(1378);
     when "010101100011" => data <= sine_rom(1379);
     when "010101100100" => data <= sine_rom(1380);
     when "010101100101" => data <= sine_rom(1381);
     when "010101100110" => data <= sine_rom(1382);
     when "010101100111" => data <= sine_rom(1383);
     when "010101101000" => data <= sine_rom(1384);
     when "010101101001" => data <= sine_rom(1385);
     when "010101101010" => data <= sine_rom(1386);
     when "010101101011" => data <= sine_rom(1387);
     when "010101101100" => data <= sine_rom(1388);
     when "010101101101" => data <= sine_rom(1389);
     when "010101101110" => data <= sine_rom(1390);
     when "010101101111" => data <= sine_rom(1391);
     when "010101110000" => data <= sine_rom(1392);
     when "010101110001" => data <= sine_rom(1393);
     when "010101110010" => data <= sine_rom(1394);
     when "010101110011" => data <= sine_rom(1395);
     when "010101110100" => data <= sine_rom(1396);
     when "010101110101" => data <= sine_rom(1397);
     when "010101110110" => data <= sine_rom(1398);
     when "010101110111" => data <= sine_rom(1399);
     when "010101111000" => data <= sine_rom(1400);
     when "010101111001" => data <= sine_rom(1401);
     when "010101111010" => data <= sine_rom(1402);
     when "010101111011" => data <= sine_rom(1403);
     when "010101111100" => data <= sine_rom(1404);
     when "010101111101" => data <= sine_rom(1405);
     when "010101111110" => data <= sine_rom(1406);
     when "010101111111" => data <= sine_rom(1407);
     when "010110000000" => data <= sine_rom(1408);
     when "010110000001" => data <= sine_rom(1409);
     when "010110000010" => data <= sine_rom(1410);
     when "010110000011" => data <= sine_rom(1411);
     when "010110000100" => data <= sine_rom(1412);
     when "010110000101" => data <= sine_rom(1413);
     when "010110000110" => data <= sine_rom(1414);
     when "010110000111" => data <= sine_rom(1415);
     when "010110001000" => data <= sine_rom(1416);
     when "010110001001" => data <= sine_rom(1417);
     when "010110001010" => data <= sine_rom(1418);
     when "010110001011" => data <= sine_rom(1419);
     when "010110001100" => data <= sine_rom(1420);
     when "010110001101" => data <= sine_rom(1421);
     when "010110001110" => data <= sine_rom(1422);
     when "010110001111" => data <= sine_rom(1423);
     when "010110010000" => data <= sine_rom(1424);
     when "010110010001" => data <= sine_rom(1425);
     when "010110010010" => data <= sine_rom(1426);
     when "010110010011" => data <= sine_rom(1427);
     when "010110010100" => data <= sine_rom(1428);
     when "010110010101" => data <= sine_rom(1429);
     when "010110010110" => data <= sine_rom(1430);
     when "010110010111" => data <= sine_rom(1431);
     when "010110011000" => data <= sine_rom(1432);
     when "010110011001" => data <= sine_rom(1433);
     when "010110011010" => data <= sine_rom(1434);
     when "010110011011" => data <= sine_rom(1435);
     when "010110011100" => data <= sine_rom(1436);
     when "010110011101" => data <= sine_rom(1437);
     when "010110011110" => data <= sine_rom(1438);
     when "010110011111" => data <= sine_rom(1439);
     when "010110100000" => data <= sine_rom(1440);
     when "010110100001" => data <= sine_rom(1441);
     when "010110100010" => data <= sine_rom(1442);
     when "010110100011" => data <= sine_rom(1443);
     when "010110100100" => data <= sine_rom(1444);
     when "010110100101" => data <= sine_rom(1445);
     when "010110100110" => data <= sine_rom(1446);
     when "010110100111" => data <= sine_rom(1447);
     when "010110101000" => data <= sine_rom(1448);
     when "010110101001" => data <= sine_rom(1449);
     when "010110101010" => data <= sine_rom(1450);
     when "010110101011" => data <= sine_rom(1451);
     when "010110101100" => data <= sine_rom(1452);
     when "010110101101" => data <= sine_rom(1453);
     when "010110101110" => data <= sine_rom(1454);
     when "010110101111" => data <= sine_rom(1455);
     when "010110110000" => data <= sine_rom(1456);
     when "010110110001" => data <= sine_rom(1457);
     when "010110110010" => data <= sine_rom(1458);
     when "010110110011" => data <= sine_rom(1459);
     when "010110110100" => data <= sine_rom(1460);
     when "010110110101" => data <= sine_rom(1461);
     when "010110110110" => data <= sine_rom(1462);
     when "010110110111" => data <= sine_rom(1463);
     when "010110111000" => data <= sine_rom(1464);
     when "010110111001" => data <= sine_rom(1465);
     when "010110111010" => data <= sine_rom(1466);
     when "010110111011" => data <= sine_rom(1467);
     when "010110111100" => data <= sine_rom(1468);
     when "010110111101" => data <= sine_rom(1469);
     when "010110111110" => data <= sine_rom(1470);
     when "010110111111" => data <= sine_rom(1471);
     when "010111000000" => data <= sine_rom(1472);
     when "010111000001" => data <= sine_rom(1473);
     when "010111000010" => data <= sine_rom(1474);
     when "010111000011" => data <= sine_rom(1475);
     when "010111000100" => data <= sine_rom(1476);
     when "010111000101" => data <= sine_rom(1477);
     when "010111000110" => data <= sine_rom(1478);
     when "010111000111" => data <= sine_rom(1479);
     when "010111001000" => data <= sine_rom(1480);
     when "010111001001" => data <= sine_rom(1481);
     when "010111001010" => data <= sine_rom(1482);
     when "010111001011" => data <= sine_rom(1483);
     when "010111001100" => data <= sine_rom(1484);
     when "010111001101" => data <= sine_rom(1485);
     when "010111001110" => data <= sine_rom(1486);
     when "010111001111" => data <= sine_rom(1487);
     when "010111010000" => data <= sine_rom(1488);
     when "010111010001" => data <= sine_rom(1489);
     when "010111010010" => data <= sine_rom(1490);
     when "010111010011" => data <= sine_rom(1491);
     when "010111010100" => data <= sine_rom(1492);
     when "010111010101" => data <= sine_rom(1493);
     when "010111010110" => data <= sine_rom(1494);
     when "010111010111" => data <= sine_rom(1495);
     when "010111011000" => data <= sine_rom(1496);
     when "010111011001" => data <= sine_rom(1497);
     when "010111011010" => data <= sine_rom(1498);
     when "010111011011" => data <= sine_rom(1499);
     when "010111011100" => data <= sine_rom(1500);
     when "010111011101" => data <= sine_rom(1501);
     when "010111011110" => data <= sine_rom(1502);
     when "010111011111" => data <= sine_rom(1503);
     when "010111100000" => data <= sine_rom(1504);
     when "010111100001" => data <= sine_rom(1505);
     when "010111100010" => data <= sine_rom(1506);
     when "010111100011" => data <= sine_rom(1507);
     when "010111100100" => data <= sine_rom(1508);
     when "010111100101" => data <= sine_rom(1509);
     when "010111100110" => data <= sine_rom(1510);
     when "010111100111" => data <= sine_rom(1511);
     when "010111101000" => data <= sine_rom(1512);
     when "010111101001" => data <= sine_rom(1513);
     when "010111101010" => data <= sine_rom(1514);
     when "010111101011" => data <= sine_rom(1515);
     when "010111101100" => data <= sine_rom(1516);
     when "010111101101" => data <= sine_rom(1517);
     when "010111101110" => data <= sine_rom(1518);
     when "010111101111" => data <= sine_rom(1519);
     when "010111110000" => data <= sine_rom(1520);
     when "010111110001" => data <= sine_rom(1521);
     when "010111110010" => data <= sine_rom(1522);
     when "010111110011" => data <= sine_rom(1523);
     when "010111110100" => data <= sine_rom(1524);
     when "010111110101" => data <= sine_rom(1525);
     when "010111110110" => data <= sine_rom(1526);
     when "010111110111" => data <= sine_rom(1527);
     when "010111111000" => data <= sine_rom(1528);
     when "010111111001" => data <= sine_rom(1529);
     when "010111111010" => data <= sine_rom(1530);
     when "010111111011" => data <= sine_rom(1531);
     when "010111111100" => data <= sine_rom(1532);
     when "010111111101" => data <= sine_rom(1533);
     when "010111111110" => data <= sine_rom(1534);
     when "010111111111" => data <= sine_rom(1535);
     when "011000000000" => data <= sine_rom(1536);
     when "011000000001" => data <= sine_rom(1537);
     when "011000000010" => data <= sine_rom(1538);
     when "011000000011" => data <= sine_rom(1539);
     when "011000000100" => data <= sine_rom(1540);
     when "011000000101" => data <= sine_rom(1541);
     when "011000000110" => data <= sine_rom(1542);
     when "011000000111" => data <= sine_rom(1543);
     when "011000001000" => data <= sine_rom(1544);
     when "011000001001" => data <= sine_rom(1545);
     when "011000001010" => data <= sine_rom(1546);
     when "011000001011" => data <= sine_rom(1547);
     when "011000001100" => data <= sine_rom(1548);
     when "011000001101" => data <= sine_rom(1549);
     when "011000001110" => data <= sine_rom(1550);
     when "011000001111" => data <= sine_rom(1551);
     when "011000010000" => data <= sine_rom(1552);
     when "011000010001" => data <= sine_rom(1553);
     when "011000010010" => data <= sine_rom(1554);
     when "011000010011" => data <= sine_rom(1555);
     when "011000010100" => data <= sine_rom(1556);
     when "011000010101" => data <= sine_rom(1557);
     when "011000010110" => data <= sine_rom(1558);
     when "011000010111" => data <= sine_rom(1559);
     when "011000011000" => data <= sine_rom(1560);
     when "011000011001" => data <= sine_rom(1561);
     when "011000011010" => data <= sine_rom(1562);
     when "011000011011" => data <= sine_rom(1563);
     when "011000011100" => data <= sine_rom(1564);
     when "011000011101" => data <= sine_rom(1565);
     when "011000011110" => data <= sine_rom(1566);
     when "011000011111" => data <= sine_rom(1567);
     when "011000100000" => data <= sine_rom(1568);
     when "011000100001" => data <= sine_rom(1569);
     when "011000100010" => data <= sine_rom(1570);
     when "011000100011" => data <= sine_rom(1571);
     when "011000100100" => data <= sine_rom(1572);
     when "011000100101" => data <= sine_rom(1573);
     when "011000100110" => data <= sine_rom(1574);
     when "011000100111" => data <= sine_rom(1575);
     when "011000101000" => data <= sine_rom(1576);
     when "011000101001" => data <= sine_rom(1577);
     when "011000101010" => data <= sine_rom(1578);
     when "011000101011" => data <= sine_rom(1579);
     when "011000101100" => data <= sine_rom(1580);
     when "011000101101" => data <= sine_rom(1581);
     when "011000101110" => data <= sine_rom(1582);
     when "011000101111" => data <= sine_rom(1583);
     when "011000110000" => data <= sine_rom(1584);
     when "011000110001" => data <= sine_rom(1585);
     when "011000110010" => data <= sine_rom(1586);
     when "011000110011" => data <= sine_rom(1587);
     when "011000110100" => data <= sine_rom(1588);
     when "011000110101" => data <= sine_rom(1589);
     when "011000110110" => data <= sine_rom(1590);
     when "011000110111" => data <= sine_rom(1591);
     when "011000111000" => data <= sine_rom(1592);
     when "011000111001" => data <= sine_rom(1593);
     when "011000111010" => data <= sine_rom(1594);
     when "011000111011" => data <= sine_rom(1595);
     when "011000111100" => data <= sine_rom(1596);
     when "011000111101" => data <= sine_rom(1597);
     when "011000111110" => data <= sine_rom(1598);
     when "011000111111" => data <= sine_rom(1599);
     when "011001000000" => data <= sine_rom(1600);
     when "011001000001" => data <= sine_rom(1601);
     when "011001000010" => data <= sine_rom(1602);
     when "011001000011" => data <= sine_rom(1603);
     when "011001000100" => data <= sine_rom(1604);
     when "011001000101" => data <= sine_rom(1605);
     when "011001000110" => data <= sine_rom(1606);
     when "011001000111" => data <= sine_rom(1607);
     when "011001001000" => data <= sine_rom(1608);
     when "011001001001" => data <= sine_rom(1609);
     when "011001001010" => data <= sine_rom(1610);
     when "011001001011" => data <= sine_rom(1611);
     when "011001001100" => data <= sine_rom(1612);
     when "011001001101" => data <= sine_rom(1613);
     when "011001001110" => data <= sine_rom(1614);
     when "011001001111" => data <= sine_rom(1615);
     when "011001010000" => data <= sine_rom(1616);
     when "011001010001" => data <= sine_rom(1617);
     when "011001010010" => data <= sine_rom(1618);
     when "011001010011" => data <= sine_rom(1619);
     when "011001010100" => data <= sine_rom(1620);
     when "011001010101" => data <= sine_rom(1621);
     when "011001010110" => data <= sine_rom(1622);
     when "011001010111" => data <= sine_rom(1623);
     when "011001011000" => data <= sine_rom(1624);
     when "011001011001" => data <= sine_rom(1625);
     when "011001011010" => data <= sine_rom(1626);
     when "011001011011" => data <= sine_rom(1627);
     when "011001011100" => data <= sine_rom(1628);
     when "011001011101" => data <= sine_rom(1629);
     when "011001011110" => data <= sine_rom(1630);
     when "011001011111" => data <= sine_rom(1631);
     when "011001100000" => data <= sine_rom(1632);
     when "011001100001" => data <= sine_rom(1633);
     when "011001100010" => data <= sine_rom(1634);
     when "011001100011" => data <= sine_rom(1635);
     when "011001100100" => data <= sine_rom(1636);
     when "011001100101" => data <= sine_rom(1637);
     when "011001100110" => data <= sine_rom(1638);
     when "011001100111" => data <= sine_rom(1639);
     when "011001101000" => data <= sine_rom(1640);
     when "011001101001" => data <= sine_rom(1641);
     when "011001101010" => data <= sine_rom(1642);
     when "011001101011" => data <= sine_rom(1643);
     when "011001101100" => data <= sine_rom(1644);
     when "011001101101" => data <= sine_rom(1645);
     when "011001101110" => data <= sine_rom(1646);
     when "011001101111" => data <= sine_rom(1647);
     when "011001110000" => data <= sine_rom(1648);
     when "011001110001" => data <= sine_rom(1649);
     when "011001110010" => data <= sine_rom(1650);
     when "011001110011" => data <= sine_rom(1651);
     when "011001110100" => data <= sine_rom(1652);
     when "011001110101" => data <= sine_rom(1653);
     when "011001110110" => data <= sine_rom(1654);
     when "011001110111" => data <= sine_rom(1655);
     when "011001111000" => data <= sine_rom(1656);
     when "011001111001" => data <= sine_rom(1657);
     when "011001111010" => data <= sine_rom(1658);
     when "011001111011" => data <= sine_rom(1659);
     when "011001111100" => data <= sine_rom(1660);
     when "011001111101" => data <= sine_rom(1661);
     when "011001111110" => data <= sine_rom(1662);
     when "011001111111" => data <= sine_rom(1663);
     when "011010000000" => data <= sine_rom(1664);
     when "011010000001" => data <= sine_rom(1665);
     when "011010000010" => data <= sine_rom(1666);
     when "011010000011" => data <= sine_rom(1667);
     when "011010000100" => data <= sine_rom(1668);
     when "011010000101" => data <= sine_rom(1669);
     when "011010000110" => data <= sine_rom(1670);
     when "011010000111" => data <= sine_rom(1671);
     when "011010001000" => data <= sine_rom(1672);
     when "011010001001" => data <= sine_rom(1673);
     when "011010001010" => data <= sine_rom(1674);
     when "011010001011" => data <= sine_rom(1675);
     when "011010001100" => data <= sine_rom(1676);
     when "011010001101" => data <= sine_rom(1677);
     when "011010001110" => data <= sine_rom(1678);
     when "011010001111" => data <= sine_rom(1679);
     when "011010010000" => data <= sine_rom(1680);
     when "011010010001" => data <= sine_rom(1681);
     when "011010010010" => data <= sine_rom(1682);
     when "011010010011" => data <= sine_rom(1683);
     when "011010010100" => data <= sine_rom(1684);
     when "011010010101" => data <= sine_rom(1685);
     when "011010010110" => data <= sine_rom(1686);
     when "011010010111" => data <= sine_rom(1687);
     when "011010011000" => data <= sine_rom(1688);
     when "011010011001" => data <= sine_rom(1689);
     when "011010011010" => data <= sine_rom(1690);
     when "011010011011" => data <= sine_rom(1691);
     when "011010011100" => data <= sine_rom(1692);
     when "011010011101" => data <= sine_rom(1693);
     when "011010011110" => data <= sine_rom(1694);
     when "011010011111" => data <= sine_rom(1695);
     when "011010100000" => data <= sine_rom(1696);
     when "011010100001" => data <= sine_rom(1697);
     when "011010100010" => data <= sine_rom(1698);
     when "011010100011" => data <= sine_rom(1699);
     when "011010100100" => data <= sine_rom(1700);
     when "011010100101" => data <= sine_rom(1701);
     when "011010100110" => data <= sine_rom(1702);
     when "011010100111" => data <= sine_rom(1703);
     when "011010101000" => data <= sine_rom(1704);
     when "011010101001" => data <= sine_rom(1705);
     when "011010101010" => data <= sine_rom(1706);
     when "011010101011" => data <= sine_rom(1707);
     when "011010101100" => data <= sine_rom(1708);
     when "011010101101" => data <= sine_rom(1709);
     when "011010101110" => data <= sine_rom(1710);
     when "011010101111" => data <= sine_rom(1711);
     when "011010110000" => data <= sine_rom(1712);
     when "011010110001" => data <= sine_rom(1713);
     when "011010110010" => data <= sine_rom(1714);
     when "011010110011" => data <= sine_rom(1715);
     when "011010110100" => data <= sine_rom(1716);
     when "011010110101" => data <= sine_rom(1717);
     when "011010110110" => data <= sine_rom(1718);
     when "011010110111" => data <= sine_rom(1719);
     when "011010111000" => data <= sine_rom(1720);
     when "011010111001" => data <= sine_rom(1721);
     when "011010111010" => data <= sine_rom(1722);
     when "011010111011" => data <= sine_rom(1723);
     when "011010111100" => data <= sine_rom(1724);
     when "011010111101" => data <= sine_rom(1725);
     when "011010111110" => data <= sine_rom(1726);
     when "011010111111" => data <= sine_rom(1727);
     when "011011000000" => data <= sine_rom(1728);
     when "011011000001" => data <= sine_rom(1729);
     when "011011000010" => data <= sine_rom(1730);
     when "011011000011" => data <= sine_rom(1731);
     when "011011000100" => data <= sine_rom(1732);
     when "011011000101" => data <= sine_rom(1733);
     when "011011000110" => data <= sine_rom(1734);
     when "011011000111" => data <= sine_rom(1735);
     when "011011001000" => data <= sine_rom(1736);
     when "011011001001" => data <= sine_rom(1737);
     when "011011001010" => data <= sine_rom(1738);
     when "011011001011" => data <= sine_rom(1739);
     when "011011001100" => data <= sine_rom(1740);
     when "011011001101" => data <= sine_rom(1741);
     when "011011001110" => data <= sine_rom(1742);
     when "011011001111" => data <= sine_rom(1743);
     when "011011010000" => data <= sine_rom(1744);
     when "011011010001" => data <= sine_rom(1745);
     when "011011010010" => data <= sine_rom(1746);
     when "011011010011" => data <= sine_rom(1747);
     when "011011010100" => data <= sine_rom(1748);
     when "011011010101" => data <= sine_rom(1749);
     when "011011010110" => data <= sine_rom(1750);
     when "011011010111" => data <= sine_rom(1751);
     when "011011011000" => data <= sine_rom(1752);
     when "011011011001" => data <= sine_rom(1753);
     when "011011011010" => data <= sine_rom(1754);
     when "011011011011" => data <= sine_rom(1755);
     when "011011011100" => data <= sine_rom(1756);
     when "011011011101" => data <= sine_rom(1757);
     when "011011011110" => data <= sine_rom(1758);
     when "011011011111" => data <= sine_rom(1759);
     when "011011100000" => data <= sine_rom(1760);
     when "011011100001" => data <= sine_rom(1761);
     when "011011100010" => data <= sine_rom(1762);
     when "011011100011" => data <= sine_rom(1763);
     when "011011100100" => data <= sine_rom(1764);
     when "011011100101" => data <= sine_rom(1765);
     when "011011100110" => data <= sine_rom(1766);
     when "011011100111" => data <= sine_rom(1767);
     when "011011101000" => data <= sine_rom(1768);
     when "011011101001" => data <= sine_rom(1769);
     when "011011101010" => data <= sine_rom(1770);
     when "011011101011" => data <= sine_rom(1771);
     when "011011101100" => data <= sine_rom(1772);
     when "011011101101" => data <= sine_rom(1773);
     when "011011101110" => data <= sine_rom(1774);
     when "011011101111" => data <= sine_rom(1775);
     when "011011110000" => data <= sine_rom(1776);
     when "011011110001" => data <= sine_rom(1777);
     when "011011110010" => data <= sine_rom(1778);
     when "011011110011" => data <= sine_rom(1779);
     when "011011110100" => data <= sine_rom(1780);
     when "011011110101" => data <= sine_rom(1781);
     when "011011110110" => data <= sine_rom(1782);
     when "011011110111" => data <= sine_rom(1783);
     when "011011111000" => data <= sine_rom(1784);
     when "011011111001" => data <= sine_rom(1785);
     when "011011111010" => data <= sine_rom(1786);
     when "011011111011" => data <= sine_rom(1787);
     when "011011111100" => data <= sine_rom(1788);
     when "011011111101" => data <= sine_rom(1789);
     when "011011111110" => data <= sine_rom(1790);
     when "011011111111" => data <= sine_rom(1791);
     when "011100000000" => data <= sine_rom(1792);
     when "011100000001" => data <= sine_rom(1793);
     when "011100000010" => data <= sine_rom(1794);
     when "011100000011" => data <= sine_rom(1795);
     when "011100000100" => data <= sine_rom(1796);
     when "011100000101" => data <= sine_rom(1797);
     when "011100000110" => data <= sine_rom(1798);
     when "011100000111" => data <= sine_rom(1799);
     when "011100001000" => data <= sine_rom(1800);
     when "011100001001" => data <= sine_rom(1801);
     when "011100001010" => data <= sine_rom(1802);
     when "011100001011" => data <= sine_rom(1803);
     when "011100001100" => data <= sine_rom(1804);
     when "011100001101" => data <= sine_rom(1805);
     when "011100001110" => data <= sine_rom(1806);
     when "011100001111" => data <= sine_rom(1807);
     when "011100010000" => data <= sine_rom(1808);
     when "011100010001" => data <= sine_rom(1809);
     when "011100010010" => data <= sine_rom(1810);
     when "011100010011" => data <= sine_rom(1811);
     when "011100010100" => data <= sine_rom(1812);
     when "011100010101" => data <= sine_rom(1813);
     when "011100010110" => data <= sine_rom(1814);
     when "011100010111" => data <= sine_rom(1815);
     when "011100011000" => data <= sine_rom(1816);
     when "011100011001" => data <= sine_rom(1817);
     when "011100011010" => data <= sine_rom(1818);
     when "011100011011" => data <= sine_rom(1819);
     when "011100011100" => data <= sine_rom(1820);
     when "011100011101" => data <= sine_rom(1821);
     when "011100011110" => data <= sine_rom(1822);
     when "011100011111" => data <= sine_rom(1823);
     when "011100100000" => data <= sine_rom(1824);
     when "011100100001" => data <= sine_rom(1825);
     when "011100100010" => data <= sine_rom(1826);
     when "011100100011" => data <= sine_rom(1827);
     when "011100100100" => data <= sine_rom(1828);
     when "011100100101" => data <= sine_rom(1829);
     when "011100100110" => data <= sine_rom(1830);
     when "011100100111" => data <= sine_rom(1831);
     when "011100101000" => data <= sine_rom(1832);
     when "011100101001" => data <= sine_rom(1833);
     when "011100101010" => data <= sine_rom(1834);
     when "011100101011" => data <= sine_rom(1835);
     when "011100101100" => data <= sine_rom(1836);
     when "011100101101" => data <= sine_rom(1837);
     when "011100101110" => data <= sine_rom(1838);
     when "011100101111" => data <= sine_rom(1839);
     when "011100110000" => data <= sine_rom(1840);
     when "011100110001" => data <= sine_rom(1841);
     when "011100110010" => data <= sine_rom(1842);
     when "011100110011" => data <= sine_rom(1843);
     when "011100110100" => data <= sine_rom(1844);
     when "011100110101" => data <= sine_rom(1845);
     when "011100110110" => data <= sine_rom(1846);
     when "011100110111" => data <= sine_rom(1847);
     when "011100111000" => data <= sine_rom(1848);
     when "011100111001" => data <= sine_rom(1849);
     when "011100111010" => data <= sine_rom(1850);
     when "011100111011" => data <= sine_rom(1851);
     when "011100111100" => data <= sine_rom(1852);
     when "011100111101" => data <= sine_rom(1853);
     when "011100111110" => data <= sine_rom(1854);
     when "011100111111" => data <= sine_rom(1855);
     when "011101000000" => data <= sine_rom(1856);
     when "011101000001" => data <= sine_rom(1857);
     when "011101000010" => data <= sine_rom(1858);
     when "011101000011" => data <= sine_rom(1859);
     when "011101000100" => data <= sine_rom(1860);
     when "011101000101" => data <= sine_rom(1861);
     when "011101000110" => data <= sine_rom(1862);
     when "011101000111" => data <= sine_rom(1863);
     when "011101001000" => data <= sine_rom(1864);
     when "011101001001" => data <= sine_rom(1865);
     when "011101001010" => data <= sine_rom(1866);
     when "011101001011" => data <= sine_rom(1867);
     when "011101001100" => data <= sine_rom(1868);
     when "011101001101" => data <= sine_rom(1869);
     when "011101001110" => data <= sine_rom(1870);
     when "011101001111" => data <= sine_rom(1871);
     when "011101010000" => data <= sine_rom(1872);
     when "011101010001" => data <= sine_rom(1873);
     when "011101010010" => data <= sine_rom(1874);
     when "011101010011" => data <= sine_rom(1875);
     when "011101010100" => data <= sine_rom(1876);
     when "011101010101" => data <= sine_rom(1877);
     when "011101010110" => data <= sine_rom(1878);
     when "011101010111" => data <= sine_rom(1879);
     when "011101011000" => data <= sine_rom(1880);
     when "011101011001" => data <= sine_rom(1881);
     when "011101011010" => data <= sine_rom(1882);
     when "011101011011" => data <= sine_rom(1883);
     when "011101011100" => data <= sine_rom(1884);
     when "011101011101" => data <= sine_rom(1885);
     when "011101011110" => data <= sine_rom(1886);
     when "011101011111" => data <= sine_rom(1887);
     when "011101100000" => data <= sine_rom(1888);
     when "011101100001" => data <= sine_rom(1889);
     when "011101100010" => data <= sine_rom(1890);
     when "011101100011" => data <= sine_rom(1891);
     when "011101100100" => data <= sine_rom(1892);
     when "011101100101" => data <= sine_rom(1893);
     when "011101100110" => data <= sine_rom(1894);
     when "011101100111" => data <= sine_rom(1895);
     when "011101101000" => data <= sine_rom(1896);
     when "011101101001" => data <= sine_rom(1897);
     when "011101101010" => data <= sine_rom(1898);
     when "011101101011" => data <= sine_rom(1899);
     when "011101101100" => data <= sine_rom(1900);
     when "011101101101" => data <= sine_rom(1901);
     when "011101101110" => data <= sine_rom(1902);
     when "011101101111" => data <= sine_rom(1903);
     when "011101110000" => data <= sine_rom(1904);
     when "011101110001" => data <= sine_rom(1905);
     when "011101110010" => data <= sine_rom(1906);
     when "011101110011" => data <= sine_rom(1907);
     when "011101110100" => data <= sine_rom(1908);
     when "011101110101" => data <= sine_rom(1909);
     when "011101110110" => data <= sine_rom(1910);
     when "011101110111" => data <= sine_rom(1911);
     when "011101111000" => data <= sine_rom(1912);
     when "011101111001" => data <= sine_rom(1913);
     when "011101111010" => data <= sine_rom(1914);
     when "011101111011" => data <= sine_rom(1915);
     when "011101111100" => data <= sine_rom(1916);
     when "011101111101" => data <= sine_rom(1917);
     when "011101111110" => data <= sine_rom(1918);
     when "011101111111" => data <= sine_rom(1919);
     when "011110000000" => data <= sine_rom(1920);
     when "011110000001" => data <= sine_rom(1921);
     when "011110000010" => data <= sine_rom(1922);
     when "011110000011" => data <= sine_rom(1923);
     when "011110000100" => data <= sine_rom(1924);
     when "011110000101" => data <= sine_rom(1925);
     when "011110000110" => data <= sine_rom(1926);
     when "011110000111" => data <= sine_rom(1927);
     when "011110001000" => data <= sine_rom(1928);
     when "011110001001" => data <= sine_rom(1929);
     when "011110001010" => data <= sine_rom(1930);
     when "011110001011" => data <= sine_rom(1931);
     when "011110001100" => data <= sine_rom(1932);
     when "011110001101" => data <= sine_rom(1933);
     when "011110001110" => data <= sine_rom(1934);
     when "011110001111" => data <= sine_rom(1935);
     when "011110010000" => data <= sine_rom(1936);
     when "011110010001" => data <= sine_rom(1937);
     when "011110010010" => data <= sine_rom(1938);
     when "011110010011" => data <= sine_rom(1939);
     when "011110010100" => data <= sine_rom(1940);
     when "011110010101" => data <= sine_rom(1941);
     when "011110010110" => data <= sine_rom(1942);
     when "011110010111" => data <= sine_rom(1943);
     when "011110011000" => data <= sine_rom(1944);
     when "011110011001" => data <= sine_rom(1945);
     when "011110011010" => data <= sine_rom(1946);
     when "011110011011" => data <= sine_rom(1947);
     when "011110011100" => data <= sine_rom(1948);
     when "011110011101" => data <= sine_rom(1949);
     when "011110011110" => data <= sine_rom(1950);
     when "011110011111" => data <= sine_rom(1951);
     when "011110100000" => data <= sine_rom(1952);
     when "011110100001" => data <= sine_rom(1953);
     when "011110100010" => data <= sine_rom(1954);
     when "011110100011" => data <= sine_rom(1955);
     when "011110100100" => data <= sine_rom(1956);
     when "011110100101" => data <= sine_rom(1957);
     when "011110100110" => data <= sine_rom(1958);
     when "011110100111" => data <= sine_rom(1959);
     when "011110101000" => data <= sine_rom(1960);
     when "011110101001" => data <= sine_rom(1961);
     when "011110101010" => data <= sine_rom(1962);
     when "011110101011" => data <= sine_rom(1963);
     when "011110101100" => data <= sine_rom(1964);
     when "011110101101" => data <= sine_rom(1965);
     when "011110101110" => data <= sine_rom(1966);
     when "011110101111" => data <= sine_rom(1967);
     when "011110110000" => data <= sine_rom(1968);
     when "011110110001" => data <= sine_rom(1969);
     when "011110110010" => data <= sine_rom(1970);
     when "011110110011" => data <= sine_rom(1971);
     when "011110110100" => data <= sine_rom(1972);
     when "011110110101" => data <= sine_rom(1973);
     when "011110110110" => data <= sine_rom(1974);
     when "011110110111" => data <= sine_rom(1975);
     when "011110111000" => data <= sine_rom(1976);
     when "011110111001" => data <= sine_rom(1977);
     when "011110111010" => data <= sine_rom(1978);
     when "011110111011" => data <= sine_rom(1979);
     when "011110111100" => data <= sine_rom(1980);
     when "011110111101" => data <= sine_rom(1981);
     when "011110111110" => data <= sine_rom(1982);
     when "011110111111" => data <= sine_rom(1983);
     when "011111000000" => data <= sine_rom(1984);
     when "011111000001" => data <= sine_rom(1985);
     when "011111000010" => data <= sine_rom(1986);
     when "011111000011" => data <= sine_rom(1987);
     when "011111000100" => data <= sine_rom(1988);
     when "011111000101" => data <= sine_rom(1989);
     when "011111000110" => data <= sine_rom(1990);
     when "011111000111" => data <= sine_rom(1991);
     when "011111001000" => data <= sine_rom(1992);
     when "011111001001" => data <= sine_rom(1993);
     when "011111001010" => data <= sine_rom(1994);
     when "011111001011" => data <= sine_rom(1995);
     when "011111001100" => data <= sine_rom(1996);
     when "011111001101" => data <= sine_rom(1997);
     when "011111001110" => data <= sine_rom(1998);
     when "011111001111" => data <= sine_rom(1999);
     when "011111010000" => data <= sine_rom(2000);
     when "011111010001" => data <= sine_rom(2001);
     when "011111010010" => data <= sine_rom(2002);
     when "011111010011" => data <= sine_rom(2003);
     when "011111010100" => data <= sine_rom(2004);
     when "011111010101" => data <= sine_rom(2005);
     when "011111010110" => data <= sine_rom(2006);
     when "011111010111" => data <= sine_rom(2007);
     when "011111011000" => data <= sine_rom(2008);
     when "011111011001" => data <= sine_rom(2009);
     when "011111011010" => data <= sine_rom(2010);
     when "011111011011" => data <= sine_rom(2011);
     when "011111011100" => data <= sine_rom(2012);
     when "011111011101" => data <= sine_rom(2013);
     when "011111011110" => data <= sine_rom(2014);
     when "011111011111" => data <= sine_rom(2015);
     when "011111100000" => data <= sine_rom(2016);
     when "011111100001" => data <= sine_rom(2017);
     when "011111100010" => data <= sine_rom(2018);
     when "011111100011" => data <= sine_rom(2019);
     when "011111100100" => data <= sine_rom(2020);
     when "011111100101" => data <= sine_rom(2021);
     when "011111100110" => data <= sine_rom(2022);
     when "011111100111" => data <= sine_rom(2023);
     when "011111101000" => data <= sine_rom(2024);
     when "011111101001" => data <= sine_rom(2025);
     when "011111101010" => data <= sine_rom(2026);
     when "011111101011" => data <= sine_rom(2027);
     when "011111101100" => data <= sine_rom(2028);
     when "011111101101" => data <= sine_rom(2029);
     when "011111101110" => data <= sine_rom(2030);
     when "011111101111" => data <= sine_rom(2031);
     when "011111110000" => data <= sine_rom(2032);
     when "011111110001" => data <= sine_rom(2033);
     when "011111110010" => data <= sine_rom(2034);
     when "011111110011" => data <= sine_rom(2035);
     when "011111110100" => data <= sine_rom(2036);
     when "011111110101" => data <= sine_rom(2037);
     when "011111110110" => data <= sine_rom(2038);
     when "011111110111" => data <= sine_rom(2039);
     when "011111111000" => data <= sine_rom(2040);
     when "011111111001" => data <= sine_rom(2041);
     when "011111111010" => data <= sine_rom(2042);
     when "011111111011" => data <= sine_rom(2043);
     when "011111111100" => data <= sine_rom(2044);
     when "011111111101" => data <= sine_rom(2045);
     when "011111111110" => data <= sine_rom(2046);
     when "011111111111" => data <= sine_rom(2047);
     when "100000000000" => data <= sine_rom(2048);
     when "100000000001" => data <= sine_rom(2049);
     when "100000000010" => data <= sine_rom(2050);
     when "100000000011" => data <= sine_rom(2051);
     when "100000000100" => data <= sine_rom(2052);
     when "100000000101" => data <= sine_rom(2053);
     when "100000000110" => data <= sine_rom(2054);
     when "100000000111" => data <= sine_rom(2055);
     when "100000001000" => data <= sine_rom(2056);
     when "100000001001" => data <= sine_rom(2057);
     when "100000001010" => data <= sine_rom(2058);
     when "100000001011" => data <= sine_rom(2059);
     when "100000001100" => data <= sine_rom(2060);
     when "100000001101" => data <= sine_rom(2061);
     when "100000001110" => data <= sine_rom(2062);
     when "100000001111" => data <= sine_rom(2063);
     when "100000010000" => data <= sine_rom(2064);
     when "100000010001" => data <= sine_rom(2065);
     when "100000010010" => data <= sine_rom(2066);
     when "100000010011" => data <= sine_rom(2067);
     when "100000010100" => data <= sine_rom(2068);
     when "100000010101" => data <= sine_rom(2069);
     when "100000010110" => data <= sine_rom(2070);
     when "100000010111" => data <= sine_rom(2071);
     when "100000011000" => data <= sine_rom(2072);
     when "100000011001" => data <= sine_rom(2073);
     when "100000011010" => data <= sine_rom(2074);
     when "100000011011" => data <= sine_rom(2075);
     when "100000011100" => data <= sine_rom(2076);
     when "100000011101" => data <= sine_rom(2077);
     when "100000011110" => data <= sine_rom(2078);
     when "100000011111" => data <= sine_rom(2079);
     when "100000100000" => data <= sine_rom(2080);
     when "100000100001" => data <= sine_rom(2081);
     when "100000100010" => data <= sine_rom(2082);
     when "100000100011" => data <= sine_rom(2083);
     when "100000100100" => data <= sine_rom(2084);
     when "100000100101" => data <= sine_rom(2085);
     when "100000100110" => data <= sine_rom(2086);
     when "100000100111" => data <= sine_rom(2087);
     when "100000101000" => data <= sine_rom(2088);
     when "100000101001" => data <= sine_rom(2089);
     when "100000101010" => data <= sine_rom(2090);
     when "100000101011" => data <= sine_rom(2091);
     when "100000101100" => data <= sine_rom(2092);
     when "100000101101" => data <= sine_rom(2093);
     when "100000101110" => data <= sine_rom(2094);
     when "100000101111" => data <= sine_rom(2095);
     when "100000110000" => data <= sine_rom(2096);
     when "100000110001" => data <= sine_rom(2097);
     when "100000110010" => data <= sine_rom(2098);
     when "100000110011" => data <= sine_rom(2099);
     when "100000110100" => data <= sine_rom(2100);
     when "100000110101" => data <= sine_rom(2101);
     when "100000110110" => data <= sine_rom(2102);
     when "100000110111" => data <= sine_rom(2103);
     when "100000111000" => data <= sine_rom(2104);
     when "100000111001" => data <= sine_rom(2105);
     when "100000111010" => data <= sine_rom(2106);
     when "100000111011" => data <= sine_rom(2107);
     when "100000111100" => data <= sine_rom(2108);
     when "100000111101" => data <= sine_rom(2109);
     when "100000111110" => data <= sine_rom(2110);
     when "100000111111" => data <= sine_rom(2111);
     when "100001000000" => data <= sine_rom(2112);
     when "100001000001" => data <= sine_rom(2113);
     when "100001000010" => data <= sine_rom(2114);
     when "100001000011" => data <= sine_rom(2115);
     when "100001000100" => data <= sine_rom(2116);
     when "100001000101" => data <= sine_rom(2117);
     when "100001000110" => data <= sine_rom(2118);
     when "100001000111" => data <= sine_rom(2119);
     when "100001001000" => data <= sine_rom(2120);
     when "100001001001" => data <= sine_rom(2121);
     when "100001001010" => data <= sine_rom(2122);
     when "100001001011" => data <= sine_rom(2123);
     when "100001001100" => data <= sine_rom(2124);
     when "100001001101" => data <= sine_rom(2125);
     when "100001001110" => data <= sine_rom(2126);
     when "100001001111" => data <= sine_rom(2127);
     when "100001010000" => data <= sine_rom(2128);
     when "100001010001" => data <= sine_rom(2129);
     when "100001010010" => data <= sine_rom(2130);
     when "100001010011" => data <= sine_rom(2131);
     when "100001010100" => data <= sine_rom(2132);
     when "100001010101" => data <= sine_rom(2133);
     when "100001010110" => data <= sine_rom(2134);
     when "100001010111" => data <= sine_rom(2135);
     when "100001011000" => data <= sine_rom(2136);
     when "100001011001" => data <= sine_rom(2137);
     when "100001011010" => data <= sine_rom(2138);
     when "100001011011" => data <= sine_rom(2139);
     when "100001011100" => data <= sine_rom(2140);
     when "100001011101" => data <= sine_rom(2141);
     when "100001011110" => data <= sine_rom(2142);
     when "100001011111" => data <= sine_rom(2143);
     when "100001100000" => data <= sine_rom(2144);
     when "100001100001" => data <= sine_rom(2145);
     when "100001100010" => data <= sine_rom(2146);
     when "100001100011" => data <= sine_rom(2147);
     when "100001100100" => data <= sine_rom(2148);
     when "100001100101" => data <= sine_rom(2149);
     when "100001100110" => data <= sine_rom(2150);
     when "100001100111" => data <= sine_rom(2151);
     when "100001101000" => data <= sine_rom(2152);
     when "100001101001" => data <= sine_rom(2153);
     when "100001101010" => data <= sine_rom(2154);
     when "100001101011" => data <= sine_rom(2155);
     when "100001101100" => data <= sine_rom(2156);
     when "100001101101" => data <= sine_rom(2157);
     when "100001101110" => data <= sine_rom(2158);
     when "100001101111" => data <= sine_rom(2159);
     when "100001110000" => data <= sine_rom(2160);
     when "100001110001" => data <= sine_rom(2161);
     when "100001110010" => data <= sine_rom(2162);
     when "100001110011" => data <= sine_rom(2163);
     when "100001110100" => data <= sine_rom(2164);
     when "100001110101" => data <= sine_rom(2165);
     when "100001110110" => data <= sine_rom(2166);
     when "100001110111" => data <= sine_rom(2167);
     when "100001111000" => data <= sine_rom(2168);
     when "100001111001" => data <= sine_rom(2169);
     when "100001111010" => data <= sine_rom(2170);
     when "100001111011" => data <= sine_rom(2171);
     when "100001111100" => data <= sine_rom(2172);
     when "100001111101" => data <= sine_rom(2173);
     when "100001111110" => data <= sine_rom(2174);
     when "100001111111" => data <= sine_rom(2175);
     when "100010000000" => data <= sine_rom(2176);
     when "100010000001" => data <= sine_rom(2177);
     when "100010000010" => data <= sine_rom(2178);
     when "100010000011" => data <= sine_rom(2179);
     when "100010000100" => data <= sine_rom(2180);
     when "100010000101" => data <= sine_rom(2181);
     when "100010000110" => data <= sine_rom(2182);
     when "100010000111" => data <= sine_rom(2183);
     when "100010001000" => data <= sine_rom(2184);
     when "100010001001" => data <= sine_rom(2185);
     when "100010001010" => data <= sine_rom(2186);
     when "100010001011" => data <= sine_rom(2187);
     when "100010001100" => data <= sine_rom(2188);
     when "100010001101" => data <= sine_rom(2189);
     when "100010001110" => data <= sine_rom(2190);
     when "100010001111" => data <= sine_rom(2191);
     when "100010010000" => data <= sine_rom(2192);
     when "100010010001" => data <= sine_rom(2193);
     when "100010010010" => data <= sine_rom(2194);
     when "100010010011" => data <= sine_rom(2195);
     when "100010010100" => data <= sine_rom(2196);
     when "100010010101" => data <= sine_rom(2197);
     when "100010010110" => data <= sine_rom(2198);
     when "100010010111" => data <= sine_rom(2199);
     when "100010011000" => data <= sine_rom(2200);
     when "100010011001" => data <= sine_rom(2201);
     when "100010011010" => data <= sine_rom(2202);
     when "100010011011" => data <= sine_rom(2203);
     when "100010011100" => data <= sine_rom(2204);
     when "100010011101" => data <= sine_rom(2205);
     when "100010011110" => data <= sine_rom(2206);
     when "100010011111" => data <= sine_rom(2207);
     when "100010100000" => data <= sine_rom(2208);
     when "100010100001" => data <= sine_rom(2209);
     when "100010100010" => data <= sine_rom(2210);
     when "100010100011" => data <= sine_rom(2211);
     when "100010100100" => data <= sine_rom(2212);
     when "100010100101" => data <= sine_rom(2213);
     when "100010100110" => data <= sine_rom(2214);
     when "100010100111" => data <= sine_rom(2215);
     when "100010101000" => data <= sine_rom(2216);
     when "100010101001" => data <= sine_rom(2217);
     when "100010101010" => data <= sine_rom(2218);
     when "100010101011" => data <= sine_rom(2219);
     when "100010101100" => data <= sine_rom(2220);
     when "100010101101" => data <= sine_rom(2221);
     when "100010101110" => data <= sine_rom(2222);
     when "100010101111" => data <= sine_rom(2223);
     when "100010110000" => data <= sine_rom(2224);
     when "100010110001" => data <= sine_rom(2225);
     when "100010110010" => data <= sine_rom(2226);
     when "100010110011" => data <= sine_rom(2227);
     when "100010110100" => data <= sine_rom(2228);
     when "100010110101" => data <= sine_rom(2229);
     when "100010110110" => data <= sine_rom(2230);
     when "100010110111" => data <= sine_rom(2231);
     when "100010111000" => data <= sine_rom(2232);
     when "100010111001" => data <= sine_rom(2233);
     when "100010111010" => data <= sine_rom(2234);
     when "100010111011" => data <= sine_rom(2235);
     when "100010111100" => data <= sine_rom(2236);
     when "100010111101" => data <= sine_rom(2237);
     when "100010111110" => data <= sine_rom(2238);
     when "100010111111" => data <= sine_rom(2239);
     when "100011000000" => data <= sine_rom(2240);
     when "100011000001" => data <= sine_rom(2241);
     when "100011000010" => data <= sine_rom(2242);
     when "100011000011" => data <= sine_rom(2243);
     when "100011000100" => data <= sine_rom(2244);
     when "100011000101" => data <= sine_rom(2245);
     when "100011000110" => data <= sine_rom(2246);
     when "100011000111" => data <= sine_rom(2247);
     when "100011001000" => data <= sine_rom(2248);
     when "100011001001" => data <= sine_rom(2249);
     when "100011001010" => data <= sine_rom(2250);
     when "100011001011" => data <= sine_rom(2251);
     when "100011001100" => data <= sine_rom(2252);
     when "100011001101" => data <= sine_rom(2253);
     when "100011001110" => data <= sine_rom(2254);
     when "100011001111" => data <= sine_rom(2255);
     when "100011010000" => data <= sine_rom(2256);
     when "100011010001" => data <= sine_rom(2257);
     when "100011010010" => data <= sine_rom(2258);
     when "100011010011" => data <= sine_rom(2259);
     when "100011010100" => data <= sine_rom(2260);
     when "100011010101" => data <= sine_rom(2261);
     when "100011010110" => data <= sine_rom(2262);
     when "100011010111" => data <= sine_rom(2263);
     when "100011011000" => data <= sine_rom(2264);
     when "100011011001" => data <= sine_rom(2265);
     when "100011011010" => data <= sine_rom(2266);
     when "100011011011" => data <= sine_rom(2267);
     when "100011011100" => data <= sine_rom(2268);
     when "100011011101" => data <= sine_rom(2269);
     when "100011011110" => data <= sine_rom(2270);
     when "100011011111" => data <= sine_rom(2271);
     when "100011100000" => data <= sine_rom(2272);
     when "100011100001" => data <= sine_rom(2273);
     when "100011100010" => data <= sine_rom(2274);
     when "100011100011" => data <= sine_rom(2275);
     when "100011100100" => data <= sine_rom(2276);
     when "100011100101" => data <= sine_rom(2277);
     when "100011100110" => data <= sine_rom(2278);
     when "100011100111" => data <= sine_rom(2279);
     when "100011101000" => data <= sine_rom(2280);
     when "100011101001" => data <= sine_rom(2281);
     when "100011101010" => data <= sine_rom(2282);
     when "100011101011" => data <= sine_rom(2283);
     when "100011101100" => data <= sine_rom(2284);
     when "100011101101" => data <= sine_rom(2285);
     when "100011101110" => data <= sine_rom(2286);
     when "100011101111" => data <= sine_rom(2287);
     when "100011110000" => data <= sine_rom(2288);
     when "100011110001" => data <= sine_rom(2289);
     when "100011110010" => data <= sine_rom(2290);
     when "100011110011" => data <= sine_rom(2291);
     when "100011110100" => data <= sine_rom(2292);
     when "100011110101" => data <= sine_rom(2293);
     when "100011110110" => data <= sine_rom(2294);
     when "100011110111" => data <= sine_rom(2295);
     when "100011111000" => data <= sine_rom(2296);
     when "100011111001" => data <= sine_rom(2297);
     when "100011111010" => data <= sine_rom(2298);
     when "100011111011" => data <= sine_rom(2299);
     when "100011111100" => data <= sine_rom(2300);
     when "100011111101" => data <= sine_rom(2301);
     when "100011111110" => data <= sine_rom(2302);
     when "100011111111" => data <= sine_rom(2303);
     when "100100000000" => data <= sine_rom(2304);
     when "100100000001" => data <= sine_rom(2305);
     when "100100000010" => data <= sine_rom(2306);
     when "100100000011" => data <= sine_rom(2307);
     when "100100000100" => data <= sine_rom(2308);
     when "100100000101" => data <= sine_rom(2309);
     when "100100000110" => data <= sine_rom(2310);
     when "100100000111" => data <= sine_rom(2311);
     when "100100001000" => data <= sine_rom(2312);
     when "100100001001" => data <= sine_rom(2313);
     when "100100001010" => data <= sine_rom(2314);
     when "100100001011" => data <= sine_rom(2315);
     when "100100001100" => data <= sine_rom(2316);
     when "100100001101" => data <= sine_rom(2317);
     when "100100001110" => data <= sine_rom(2318);
     when "100100001111" => data <= sine_rom(2319);
     when "100100010000" => data <= sine_rom(2320);
     when "100100010001" => data <= sine_rom(2321);
     when "100100010010" => data <= sine_rom(2322);
     when "100100010011" => data <= sine_rom(2323);
     when "100100010100" => data <= sine_rom(2324);
     when "100100010101" => data <= sine_rom(2325);
     when "100100010110" => data <= sine_rom(2326);
     when "100100010111" => data <= sine_rom(2327);
     when "100100011000" => data <= sine_rom(2328);
     when "100100011001" => data <= sine_rom(2329);
     when "100100011010" => data <= sine_rom(2330);
     when "100100011011" => data <= sine_rom(2331);
     when "100100011100" => data <= sine_rom(2332);
     when "100100011101" => data <= sine_rom(2333);
     when "100100011110" => data <= sine_rom(2334);
     when "100100011111" => data <= sine_rom(2335);
     when "100100100000" => data <= sine_rom(2336);
     when "100100100001" => data <= sine_rom(2337);
     when "100100100010" => data <= sine_rom(2338);
     when "100100100011" => data <= sine_rom(2339);
     when "100100100100" => data <= sine_rom(2340);
     when "100100100101" => data <= sine_rom(2341);
     when "100100100110" => data <= sine_rom(2342);
     when "100100100111" => data <= sine_rom(2343);
     when "100100101000" => data <= sine_rom(2344);
     when "100100101001" => data <= sine_rom(2345);
     when "100100101010" => data <= sine_rom(2346);
     when "100100101011" => data <= sine_rom(2347);
     when "100100101100" => data <= sine_rom(2348);
     when "100100101101" => data <= sine_rom(2349);
     when "100100101110" => data <= sine_rom(2350);
     when "100100101111" => data <= sine_rom(2351);
     when "100100110000" => data <= sine_rom(2352);
     when "100100110001" => data <= sine_rom(2353);
     when "100100110010" => data <= sine_rom(2354);
     when "100100110011" => data <= sine_rom(2355);
     when "100100110100" => data <= sine_rom(2356);
     when "100100110101" => data <= sine_rom(2357);
     when "100100110110" => data <= sine_rom(2358);
     when "100100110111" => data <= sine_rom(2359);
     when "100100111000" => data <= sine_rom(2360);
     when "100100111001" => data <= sine_rom(2361);
     when "100100111010" => data <= sine_rom(2362);
     when "100100111011" => data <= sine_rom(2363);
     when "100100111100" => data <= sine_rom(2364);
     when "100100111101" => data <= sine_rom(2365);
     when "100100111110" => data <= sine_rom(2366);
     when "100100111111" => data <= sine_rom(2367);
     when "100101000000" => data <= sine_rom(2368);
     when "100101000001" => data <= sine_rom(2369);
     when "100101000010" => data <= sine_rom(2370);
     when "100101000011" => data <= sine_rom(2371);
     when "100101000100" => data <= sine_rom(2372);
     when "100101000101" => data <= sine_rom(2373);
     when "100101000110" => data <= sine_rom(2374);
     when "100101000111" => data <= sine_rom(2375);
     when "100101001000" => data <= sine_rom(2376);
     when "100101001001" => data <= sine_rom(2377);
     when "100101001010" => data <= sine_rom(2378);
     when "100101001011" => data <= sine_rom(2379);
     when "100101001100" => data <= sine_rom(2380);
     when "100101001101" => data <= sine_rom(2381);
     when "100101001110" => data <= sine_rom(2382);
     when "100101001111" => data <= sine_rom(2383);
     when "100101010000" => data <= sine_rom(2384);
     when "100101010001" => data <= sine_rom(2385);
     when "100101010010" => data <= sine_rom(2386);
     when "100101010011" => data <= sine_rom(2387);
     when "100101010100" => data <= sine_rom(2388);
     when "100101010101" => data <= sine_rom(2389);
     when "100101010110" => data <= sine_rom(2390);
     when "100101010111" => data <= sine_rom(2391);
     when "100101011000" => data <= sine_rom(2392);
     when "100101011001" => data <= sine_rom(2393);
     when "100101011010" => data <= sine_rom(2394);
     when "100101011011" => data <= sine_rom(2395);
     when "100101011100" => data <= sine_rom(2396);
     when "100101011101" => data <= sine_rom(2397);
     when "100101011110" => data <= sine_rom(2398);
     when "100101011111" => data <= sine_rom(2399);
     when "100101100000" => data <= sine_rom(2400);
     when "100101100001" => data <= sine_rom(2401);
     when "100101100010" => data <= sine_rom(2402);
     when "100101100011" => data <= sine_rom(2403);
     when "100101100100" => data <= sine_rom(2404);
     when "100101100101" => data <= sine_rom(2405);
     when "100101100110" => data <= sine_rom(2406);
     when "100101100111" => data <= sine_rom(2407);
     when "100101101000" => data <= sine_rom(2408);
     when "100101101001" => data <= sine_rom(2409);
     when "100101101010" => data <= sine_rom(2410);
     when "100101101011" => data <= sine_rom(2411);
     when "100101101100" => data <= sine_rom(2412);
     when "100101101101" => data <= sine_rom(2413);
     when "100101101110" => data <= sine_rom(2414);
     when "100101101111" => data <= sine_rom(2415);
     when "100101110000" => data <= sine_rom(2416);
     when "100101110001" => data <= sine_rom(2417);
     when "100101110010" => data <= sine_rom(2418);
     when "100101110011" => data <= sine_rom(2419);
     when "100101110100" => data <= sine_rom(2420);
     when "100101110101" => data <= sine_rom(2421);
     when "100101110110" => data <= sine_rom(2422);
     when "100101110111" => data <= sine_rom(2423);
     when "100101111000" => data <= sine_rom(2424);
     when "100101111001" => data <= sine_rom(2425);
     when "100101111010" => data <= sine_rom(2426);
     when "100101111011" => data <= sine_rom(2427);
     when "100101111100" => data <= sine_rom(2428);
     when "100101111101" => data <= sine_rom(2429);
     when "100101111110" => data <= sine_rom(2430);
     when "100101111111" => data <= sine_rom(2431);
     when "100110000000" => data <= sine_rom(2432);
     when "100110000001" => data <= sine_rom(2433);
     when "100110000010" => data <= sine_rom(2434);
     when "100110000011" => data <= sine_rom(2435);
     when "100110000100" => data <= sine_rom(2436);
     when "100110000101" => data <= sine_rom(2437);
     when "100110000110" => data <= sine_rom(2438);
     when "100110000111" => data <= sine_rom(2439);
     when "100110001000" => data <= sine_rom(2440);
     when "100110001001" => data <= sine_rom(2441);
     when "100110001010" => data <= sine_rom(2442);
     when "100110001011" => data <= sine_rom(2443);
     when "100110001100" => data <= sine_rom(2444);
     when "100110001101" => data <= sine_rom(2445);
     when "100110001110" => data <= sine_rom(2446);
     when "100110001111" => data <= sine_rom(2447);
     when "100110010000" => data <= sine_rom(2448);
     when "100110010001" => data <= sine_rom(2449);
     when "100110010010" => data <= sine_rom(2450);
     when "100110010011" => data <= sine_rom(2451);
     when "100110010100" => data <= sine_rom(2452);
     when "100110010101" => data <= sine_rom(2453);
     when "100110010110" => data <= sine_rom(2454);
     when "100110010111" => data <= sine_rom(2455);
     when "100110011000" => data <= sine_rom(2456);
     when "100110011001" => data <= sine_rom(2457);
     when "100110011010" => data <= sine_rom(2458);
     when "100110011011" => data <= sine_rom(2459);
     when "100110011100" => data <= sine_rom(2460);
     when "100110011101" => data <= sine_rom(2461);
     when "100110011110" => data <= sine_rom(2462);
     when "100110011111" => data <= sine_rom(2463);
     when "100110100000" => data <= sine_rom(2464);
     when "100110100001" => data <= sine_rom(2465);
     when "100110100010" => data <= sine_rom(2466);
     when "100110100011" => data <= sine_rom(2467);
     when "100110100100" => data <= sine_rom(2468);
     when "100110100101" => data <= sine_rom(2469);
     when "100110100110" => data <= sine_rom(2470);
     when "100110100111" => data <= sine_rom(2471);
     when "100110101000" => data <= sine_rom(2472);
     when "100110101001" => data <= sine_rom(2473);
     when "100110101010" => data <= sine_rom(2474);
     when "100110101011" => data <= sine_rom(2475);
     when "100110101100" => data <= sine_rom(2476);
     when "100110101101" => data <= sine_rom(2477);
     when "100110101110" => data <= sine_rom(2478);
     when "100110101111" => data <= sine_rom(2479);
     when "100110110000" => data <= sine_rom(2480);
     when "100110110001" => data <= sine_rom(2481);
     when "100110110010" => data <= sine_rom(2482);
     when "100110110011" => data <= sine_rom(2483);
     when "100110110100" => data <= sine_rom(2484);
     when "100110110101" => data <= sine_rom(2485);
     when "100110110110" => data <= sine_rom(2486);
     when "100110110111" => data <= sine_rom(2487);
     when "100110111000" => data <= sine_rom(2488);
     when "100110111001" => data <= sine_rom(2489);
     when "100110111010" => data <= sine_rom(2490);
     when "100110111011" => data <= sine_rom(2491);
     when "100110111100" => data <= sine_rom(2492);
     when "100110111101" => data <= sine_rom(2493);
     when "100110111110" => data <= sine_rom(2494);
     when "100110111111" => data <= sine_rom(2495);
     when "100111000000" => data <= sine_rom(2496);
     when "100111000001" => data <= sine_rom(2497);
     when "100111000010" => data <= sine_rom(2498);
     when "100111000011" => data <= sine_rom(2499);
     when "100111000100" => data <= sine_rom(2500);
     when "100111000101" => data <= sine_rom(2501);
     when "100111000110" => data <= sine_rom(2502);
     when "100111000111" => data <= sine_rom(2503);
     when "100111001000" => data <= sine_rom(2504);
     when "100111001001" => data <= sine_rom(2505);
     when "100111001010" => data <= sine_rom(2506);
     when "100111001011" => data <= sine_rom(2507);
     when "100111001100" => data <= sine_rom(2508);
     when "100111001101" => data <= sine_rom(2509);
     when "100111001110" => data <= sine_rom(2510);
     when "100111001111" => data <= sine_rom(2511);
     when "100111010000" => data <= sine_rom(2512);
     when "100111010001" => data <= sine_rom(2513);
     when "100111010010" => data <= sine_rom(2514);
     when "100111010011" => data <= sine_rom(2515);
     when "100111010100" => data <= sine_rom(2516);
     when "100111010101" => data <= sine_rom(2517);
     when "100111010110" => data <= sine_rom(2518);
     when "100111010111" => data <= sine_rom(2519);
     when "100111011000" => data <= sine_rom(2520);
     when "100111011001" => data <= sine_rom(2521);
     when "100111011010" => data <= sine_rom(2522);
     when "100111011011" => data <= sine_rom(2523);
     when "100111011100" => data <= sine_rom(2524);
     when "100111011101" => data <= sine_rom(2525);
     when "100111011110" => data <= sine_rom(2526);
     when "100111011111" => data <= sine_rom(2527);
     when "100111100000" => data <= sine_rom(2528);
     when "100111100001" => data <= sine_rom(2529);
     when "100111100010" => data <= sine_rom(2530);
     when "100111100011" => data <= sine_rom(2531);
     when "100111100100" => data <= sine_rom(2532);
     when "100111100101" => data <= sine_rom(2533);
     when "100111100110" => data <= sine_rom(2534);
     when "100111100111" => data <= sine_rom(2535);
     when "100111101000" => data <= sine_rom(2536);
     when "100111101001" => data <= sine_rom(2537);
     when "100111101010" => data <= sine_rom(2538);
     when "100111101011" => data <= sine_rom(2539);
     when "100111101100" => data <= sine_rom(2540);
     when "100111101101" => data <= sine_rom(2541);
     when "100111101110" => data <= sine_rom(2542);
     when "100111101111" => data <= sine_rom(2543);
     when "100111110000" => data <= sine_rom(2544);
     when "100111110001" => data <= sine_rom(2545);
     when "100111110010" => data <= sine_rom(2546);
     when "100111110011" => data <= sine_rom(2547);
     when "100111110100" => data <= sine_rom(2548);
     when "100111110101" => data <= sine_rom(2549);
     when "100111110110" => data <= sine_rom(2550);
     when "100111110111" => data <= sine_rom(2551);
     when "100111111000" => data <= sine_rom(2552);
     when "100111111001" => data <= sine_rom(2553);
     when "100111111010" => data <= sine_rom(2554);
     when "100111111011" => data <= sine_rom(2555);
     when "100111111100" => data <= sine_rom(2556);
     when "100111111101" => data <= sine_rom(2557);
     when "100111111110" => data <= sine_rom(2558);
     when "100111111111" => data <= sine_rom(2559);
     when "101000000000" => data <= sine_rom(2560);
     when "101000000001" => data <= sine_rom(2561);
     when "101000000010" => data <= sine_rom(2562);
     when "101000000011" => data <= sine_rom(2563);
     when "101000000100" => data <= sine_rom(2564);
     when "101000000101" => data <= sine_rom(2565);
     when "101000000110" => data <= sine_rom(2566);
     when "101000000111" => data <= sine_rom(2567);
     when "101000001000" => data <= sine_rom(2568);
     when "101000001001" => data <= sine_rom(2569);
     when "101000001010" => data <= sine_rom(2570);
     when "101000001011" => data <= sine_rom(2571);
     when "101000001100" => data <= sine_rom(2572);
     when "101000001101" => data <= sine_rom(2573);
     when "101000001110" => data <= sine_rom(2574);
     when "101000001111" => data <= sine_rom(2575);
     when "101000010000" => data <= sine_rom(2576);
     when "101000010001" => data <= sine_rom(2577);
     when "101000010010" => data <= sine_rom(2578);
     when "101000010011" => data <= sine_rom(2579);
     when "101000010100" => data <= sine_rom(2580);
     when "101000010101" => data <= sine_rom(2581);
     when "101000010110" => data <= sine_rom(2582);
     when "101000010111" => data <= sine_rom(2583);
     when "101000011000" => data <= sine_rom(2584);
     when "101000011001" => data <= sine_rom(2585);
     when "101000011010" => data <= sine_rom(2586);
     when "101000011011" => data <= sine_rom(2587);
     when "101000011100" => data <= sine_rom(2588);
     when "101000011101" => data <= sine_rom(2589);
     when "101000011110" => data <= sine_rom(2590);
     when "101000011111" => data <= sine_rom(2591);
     when "101000100000" => data <= sine_rom(2592);
     when "101000100001" => data <= sine_rom(2593);
     when "101000100010" => data <= sine_rom(2594);
     when "101000100011" => data <= sine_rom(2595);
     when "101000100100" => data <= sine_rom(2596);
     when "101000100101" => data <= sine_rom(2597);
     when "101000100110" => data <= sine_rom(2598);
     when "101000100111" => data <= sine_rom(2599);
     when "101000101000" => data <= sine_rom(2600);
     when "101000101001" => data <= sine_rom(2601);
     when "101000101010" => data <= sine_rom(2602);
     when "101000101011" => data <= sine_rom(2603);
     when "101000101100" => data <= sine_rom(2604);
     when "101000101101" => data <= sine_rom(2605);
     when "101000101110" => data <= sine_rom(2606);
     when "101000101111" => data <= sine_rom(2607);
     when "101000110000" => data <= sine_rom(2608);
     when "101000110001" => data <= sine_rom(2609);
     when "101000110010" => data <= sine_rom(2610);
     when "101000110011" => data <= sine_rom(2611);
     when "101000110100" => data <= sine_rom(2612);
     when "101000110101" => data <= sine_rom(2613);
     when "101000110110" => data <= sine_rom(2614);
     when "101000110111" => data <= sine_rom(2615);
     when "101000111000" => data <= sine_rom(2616);
     when "101000111001" => data <= sine_rom(2617);
     when "101000111010" => data <= sine_rom(2618);
     when "101000111011" => data <= sine_rom(2619);
     when "101000111100" => data <= sine_rom(2620);
     when "101000111101" => data <= sine_rom(2621);
     when "101000111110" => data <= sine_rom(2622);
     when "101000111111" => data <= sine_rom(2623);
     when "101001000000" => data <= sine_rom(2624);
     when "101001000001" => data <= sine_rom(2625);
     when "101001000010" => data <= sine_rom(2626);
     when "101001000011" => data <= sine_rom(2627);
     when "101001000100" => data <= sine_rom(2628);
     when "101001000101" => data <= sine_rom(2629);
     when "101001000110" => data <= sine_rom(2630);
     when "101001000111" => data <= sine_rom(2631);
     when "101001001000" => data <= sine_rom(2632);
     when "101001001001" => data <= sine_rom(2633);
     when "101001001010" => data <= sine_rom(2634);
     when "101001001011" => data <= sine_rom(2635);
     when "101001001100" => data <= sine_rom(2636);
     when "101001001101" => data <= sine_rom(2637);
     when "101001001110" => data <= sine_rom(2638);
     when "101001001111" => data <= sine_rom(2639);
     when "101001010000" => data <= sine_rom(2640);
     when "101001010001" => data <= sine_rom(2641);
     when "101001010010" => data <= sine_rom(2642);
     when "101001010011" => data <= sine_rom(2643);
     when "101001010100" => data <= sine_rom(2644);
     when "101001010101" => data <= sine_rom(2645);
     when "101001010110" => data <= sine_rom(2646);
     when "101001010111" => data <= sine_rom(2647);
     when "101001011000" => data <= sine_rom(2648);
     when "101001011001" => data <= sine_rom(2649);
     when "101001011010" => data <= sine_rom(2650);
     when "101001011011" => data <= sine_rom(2651);
     when "101001011100" => data <= sine_rom(2652);
     when "101001011101" => data <= sine_rom(2653);
     when "101001011110" => data <= sine_rom(2654);
     when "101001011111" => data <= sine_rom(2655);
     when "101001100000" => data <= sine_rom(2656);
     when "101001100001" => data <= sine_rom(2657);
     when "101001100010" => data <= sine_rom(2658);
     when "101001100011" => data <= sine_rom(2659);
     when "101001100100" => data <= sine_rom(2660);
     when "101001100101" => data <= sine_rom(2661);
     when "101001100110" => data <= sine_rom(2662);
     when "101001100111" => data <= sine_rom(2663);
     when "101001101000" => data <= sine_rom(2664);
     when "101001101001" => data <= sine_rom(2665);
     when "101001101010" => data <= sine_rom(2666);
     when "101001101011" => data <= sine_rom(2667);
     when "101001101100" => data <= sine_rom(2668);
     when "101001101101" => data <= sine_rom(2669);
     when "101001101110" => data <= sine_rom(2670);
     when "101001101111" => data <= sine_rom(2671);
     when "101001110000" => data <= sine_rom(2672);
     when "101001110001" => data <= sine_rom(2673);
     when "101001110010" => data <= sine_rom(2674);
     when "101001110011" => data <= sine_rom(2675);
     when "101001110100" => data <= sine_rom(2676);
     when "101001110101" => data <= sine_rom(2677);
     when "101001110110" => data <= sine_rom(2678);
     when "101001110111" => data <= sine_rom(2679);
     when "101001111000" => data <= sine_rom(2680);
     when "101001111001" => data <= sine_rom(2681);
     when "101001111010" => data <= sine_rom(2682);
     when "101001111011" => data <= sine_rom(2683);
     when "101001111100" => data <= sine_rom(2684);
     when "101001111101" => data <= sine_rom(2685);
     when "101001111110" => data <= sine_rom(2686);
     when "101001111111" => data <= sine_rom(2687);
     when "101010000000" => data <= sine_rom(2688);
     when "101010000001" => data <= sine_rom(2689);
     when "101010000010" => data <= sine_rom(2690);
     when "101010000011" => data <= sine_rom(2691);
     when "101010000100" => data <= sine_rom(2692);
     when "101010000101" => data <= sine_rom(2693);
     when "101010000110" => data <= sine_rom(2694);
     when "101010000111" => data <= sine_rom(2695);
     when "101010001000" => data <= sine_rom(2696);
     when "101010001001" => data <= sine_rom(2697);
     when "101010001010" => data <= sine_rom(2698);
     when "101010001011" => data <= sine_rom(2699);
     when "101010001100" => data <= sine_rom(2700);
     when "101010001101" => data <= sine_rom(2701);
     when "101010001110" => data <= sine_rom(2702);
     when "101010001111" => data <= sine_rom(2703);
     when "101010010000" => data <= sine_rom(2704);
     when "101010010001" => data <= sine_rom(2705);
     when "101010010010" => data <= sine_rom(2706);
     when "101010010011" => data <= sine_rom(2707);
     when "101010010100" => data <= sine_rom(2708);
     when "101010010101" => data <= sine_rom(2709);
     when "101010010110" => data <= sine_rom(2710);
     when "101010010111" => data <= sine_rom(2711);
     when "101010011000" => data <= sine_rom(2712);
     when "101010011001" => data <= sine_rom(2713);
     when "101010011010" => data <= sine_rom(2714);
     when "101010011011" => data <= sine_rom(2715);
     when "101010011100" => data <= sine_rom(2716);
     when "101010011101" => data <= sine_rom(2717);
     when "101010011110" => data <= sine_rom(2718);
     when "101010011111" => data <= sine_rom(2719);
     when "101010100000" => data <= sine_rom(2720);
     when "101010100001" => data <= sine_rom(2721);
     when "101010100010" => data <= sine_rom(2722);
     when "101010100011" => data <= sine_rom(2723);
     when "101010100100" => data <= sine_rom(2724);
     when "101010100101" => data <= sine_rom(2725);
     when "101010100110" => data <= sine_rom(2726);
     when "101010100111" => data <= sine_rom(2727);
     when "101010101000" => data <= sine_rom(2728);
     when "101010101001" => data <= sine_rom(2729);
     when "101010101010" => data <= sine_rom(2730);
     when "101010101011" => data <= sine_rom(2731);
     when "101010101100" => data <= sine_rom(2732);
     when "101010101101" => data <= sine_rom(2733);
     when "101010101110" => data <= sine_rom(2734);
     when "101010101111" => data <= sine_rom(2735);
     when "101010110000" => data <= sine_rom(2736);
     when "101010110001" => data <= sine_rom(2737);
     when "101010110010" => data <= sine_rom(2738);
     when "101010110011" => data <= sine_rom(2739);
     when "101010110100" => data <= sine_rom(2740);
     when "101010110101" => data <= sine_rom(2741);
     when "101010110110" => data <= sine_rom(2742);
     when "101010110111" => data <= sine_rom(2743);
     when "101010111000" => data <= sine_rom(2744);
     when "101010111001" => data <= sine_rom(2745);
     when "101010111010" => data <= sine_rom(2746);
     when "101010111011" => data <= sine_rom(2747);
     when "101010111100" => data <= sine_rom(2748);
     when "101010111101" => data <= sine_rom(2749);
     when "101010111110" => data <= sine_rom(2750);
     when "101010111111" => data <= sine_rom(2751);
     when "101011000000" => data <= sine_rom(2752);
     when "101011000001" => data <= sine_rom(2753);
     when "101011000010" => data <= sine_rom(2754);
     when "101011000011" => data <= sine_rom(2755);
     when "101011000100" => data <= sine_rom(2756);
     when "101011000101" => data <= sine_rom(2757);
     when "101011000110" => data <= sine_rom(2758);
     when "101011000111" => data <= sine_rom(2759);
     when "101011001000" => data <= sine_rom(2760);
     when "101011001001" => data <= sine_rom(2761);
     when "101011001010" => data <= sine_rom(2762);
     when "101011001011" => data <= sine_rom(2763);
     when "101011001100" => data <= sine_rom(2764);
     when "101011001101" => data <= sine_rom(2765);
     when "101011001110" => data <= sine_rom(2766);
     when "101011001111" => data <= sine_rom(2767);
     when "101011010000" => data <= sine_rom(2768);
     when "101011010001" => data <= sine_rom(2769);
     when "101011010010" => data <= sine_rom(2770);
     when "101011010011" => data <= sine_rom(2771);
     when "101011010100" => data <= sine_rom(2772);
     when "101011010101" => data <= sine_rom(2773);
     when "101011010110" => data <= sine_rom(2774);
     when "101011010111" => data <= sine_rom(2775);
     when "101011011000" => data <= sine_rom(2776);
     when "101011011001" => data <= sine_rom(2777);
     when "101011011010" => data <= sine_rom(2778);
     when "101011011011" => data <= sine_rom(2779);
     when "101011011100" => data <= sine_rom(2780);
     when "101011011101" => data <= sine_rom(2781);
     when "101011011110" => data <= sine_rom(2782);
     when "101011011111" => data <= sine_rom(2783);
     when "101011100000" => data <= sine_rom(2784);
     when "101011100001" => data <= sine_rom(2785);
     when "101011100010" => data <= sine_rom(2786);
     when "101011100011" => data <= sine_rom(2787);
     when "101011100100" => data <= sine_rom(2788);
     when "101011100101" => data <= sine_rom(2789);
     when "101011100110" => data <= sine_rom(2790);
     when "101011100111" => data <= sine_rom(2791);
     when "101011101000" => data <= sine_rom(2792);
     when "101011101001" => data <= sine_rom(2793);
     when "101011101010" => data <= sine_rom(2794);
     when "101011101011" => data <= sine_rom(2795);
     when "101011101100" => data <= sine_rom(2796);
     when "101011101101" => data <= sine_rom(2797);
     when "101011101110" => data <= sine_rom(2798);
     when "101011101111" => data <= sine_rom(2799);
     when "101011110000" => data <= sine_rom(2800);
     when "101011110001" => data <= sine_rom(2801);
     when "101011110010" => data <= sine_rom(2802);
     when "101011110011" => data <= sine_rom(2803);
     when "101011110100" => data <= sine_rom(2804);
     when "101011110101" => data <= sine_rom(2805);
     when "101011110110" => data <= sine_rom(2806);
     when "101011110111" => data <= sine_rom(2807);
     when "101011111000" => data <= sine_rom(2808);
     when "101011111001" => data <= sine_rom(2809);
     when "101011111010" => data <= sine_rom(2810);
     when "101011111011" => data <= sine_rom(2811);
     when "101011111100" => data <= sine_rom(2812);
     when "101011111101" => data <= sine_rom(2813);
     when "101011111110" => data <= sine_rom(2814);
     when "101011111111" => data <= sine_rom(2815);
     when "101100000000" => data <= sine_rom(2816);
     when "101100000001" => data <= sine_rom(2817);
     when "101100000010" => data <= sine_rom(2818);
     when "101100000011" => data <= sine_rom(2819);
     when "101100000100" => data <= sine_rom(2820);
     when "101100000101" => data <= sine_rom(2821);
     when "101100000110" => data <= sine_rom(2822);
     when "101100000111" => data <= sine_rom(2823);
     when "101100001000" => data <= sine_rom(2824);
     when "101100001001" => data <= sine_rom(2825);
     when "101100001010" => data <= sine_rom(2826);
     when "101100001011" => data <= sine_rom(2827);
     when "101100001100" => data <= sine_rom(2828);
     when "101100001101" => data <= sine_rom(2829);
     when "101100001110" => data <= sine_rom(2830);
     when "101100001111" => data <= sine_rom(2831);
     when "101100010000" => data <= sine_rom(2832);
     when "101100010001" => data <= sine_rom(2833);
     when "101100010010" => data <= sine_rom(2834);
     when "101100010011" => data <= sine_rom(2835);
     when "101100010100" => data <= sine_rom(2836);
     when "101100010101" => data <= sine_rom(2837);
     when "101100010110" => data <= sine_rom(2838);
     when "101100010111" => data <= sine_rom(2839);
     when "101100011000" => data <= sine_rom(2840);
     when "101100011001" => data <= sine_rom(2841);
     when "101100011010" => data <= sine_rom(2842);
     when "101100011011" => data <= sine_rom(2843);
     when "101100011100" => data <= sine_rom(2844);
     when "101100011101" => data <= sine_rom(2845);
     when "101100011110" => data <= sine_rom(2846);
     when "101100011111" => data <= sine_rom(2847);
     when "101100100000" => data <= sine_rom(2848);
     when "101100100001" => data <= sine_rom(2849);
     when "101100100010" => data <= sine_rom(2850);
     when "101100100011" => data <= sine_rom(2851);
     when "101100100100" => data <= sine_rom(2852);
     when "101100100101" => data <= sine_rom(2853);
     when "101100100110" => data <= sine_rom(2854);
     when "101100100111" => data <= sine_rom(2855);
     when "101100101000" => data <= sine_rom(2856);
     when "101100101001" => data <= sine_rom(2857);
     when "101100101010" => data <= sine_rom(2858);
     when "101100101011" => data <= sine_rom(2859);
     when "101100101100" => data <= sine_rom(2860);
     when "101100101101" => data <= sine_rom(2861);
     when "101100101110" => data <= sine_rom(2862);
     when "101100101111" => data <= sine_rom(2863);
     when "101100110000" => data <= sine_rom(2864);
     when "101100110001" => data <= sine_rom(2865);
     when "101100110010" => data <= sine_rom(2866);
     when "101100110011" => data <= sine_rom(2867);
     when "101100110100" => data <= sine_rom(2868);
     when "101100110101" => data <= sine_rom(2869);
     when "101100110110" => data <= sine_rom(2870);
     when "101100110111" => data <= sine_rom(2871);
     when "101100111000" => data <= sine_rom(2872);
     when "101100111001" => data <= sine_rom(2873);
     when "101100111010" => data <= sine_rom(2874);
     when "101100111011" => data <= sine_rom(2875);
     when "101100111100" => data <= sine_rom(2876);
     when "101100111101" => data <= sine_rom(2877);
     when "101100111110" => data <= sine_rom(2878);
     when "101100111111" => data <= sine_rom(2879);
     when "101101000000" => data <= sine_rom(2880);
     when "101101000001" => data <= sine_rom(2881);
     when "101101000010" => data <= sine_rom(2882);
     when "101101000011" => data <= sine_rom(2883);
     when "101101000100" => data <= sine_rom(2884);
     when "101101000101" => data <= sine_rom(2885);
     when "101101000110" => data <= sine_rom(2886);
     when "101101000111" => data <= sine_rom(2887);
     when "101101001000" => data <= sine_rom(2888);
     when "101101001001" => data <= sine_rom(2889);
     when "101101001010" => data <= sine_rom(2890);
     when "101101001011" => data <= sine_rom(2891);
     when "101101001100" => data <= sine_rom(2892);
     when "101101001101" => data <= sine_rom(2893);
     when "101101001110" => data <= sine_rom(2894);
     when "101101001111" => data <= sine_rom(2895);
     when "101101010000" => data <= sine_rom(2896);
     when "101101010001" => data <= sine_rom(2897);
     when "101101010010" => data <= sine_rom(2898);
     when "101101010011" => data <= sine_rom(2899);
     when "101101010100" => data <= sine_rom(2900);
     when "101101010101" => data <= sine_rom(2901);
     when "101101010110" => data <= sine_rom(2902);
     when "101101010111" => data <= sine_rom(2903);
     when "101101011000" => data <= sine_rom(2904);
     when "101101011001" => data <= sine_rom(2905);
     when "101101011010" => data <= sine_rom(2906);
     when "101101011011" => data <= sine_rom(2907);
     when "101101011100" => data <= sine_rom(2908);
     when "101101011101" => data <= sine_rom(2909);
     when "101101011110" => data <= sine_rom(2910);
     when "101101011111" => data <= sine_rom(2911);
     when "101101100000" => data <= sine_rom(2912);
     when "101101100001" => data <= sine_rom(2913);
     when "101101100010" => data <= sine_rom(2914);
     when "101101100011" => data <= sine_rom(2915);
     when "101101100100" => data <= sine_rom(2916);
     when "101101100101" => data <= sine_rom(2917);
     when "101101100110" => data <= sine_rom(2918);
     when "101101100111" => data <= sine_rom(2919);
     when "101101101000" => data <= sine_rom(2920);
     when "101101101001" => data <= sine_rom(2921);
     when "101101101010" => data <= sine_rom(2922);
     when "101101101011" => data <= sine_rom(2923);
     when "101101101100" => data <= sine_rom(2924);
     when "101101101101" => data <= sine_rom(2925);
     when "101101101110" => data <= sine_rom(2926);
     when "101101101111" => data <= sine_rom(2927);
     when "101101110000" => data <= sine_rom(2928);
     when "101101110001" => data <= sine_rom(2929);
     when "101101110010" => data <= sine_rom(2930);
     when "101101110011" => data <= sine_rom(2931);
     when "101101110100" => data <= sine_rom(2932);
     when "101101110101" => data <= sine_rom(2933);
     when "101101110110" => data <= sine_rom(2934);
     when "101101110111" => data <= sine_rom(2935);
     when "101101111000" => data <= sine_rom(2936);
     when "101101111001" => data <= sine_rom(2937);
     when "101101111010" => data <= sine_rom(2938);
     when "101101111011" => data <= sine_rom(2939);
     when "101101111100" => data <= sine_rom(2940);
     when "101101111101" => data <= sine_rom(2941);
     when "101101111110" => data <= sine_rom(2942);
     when "101101111111" => data <= sine_rom(2943);
     when "101110000000" => data <= sine_rom(2944);
     when "101110000001" => data <= sine_rom(2945);
     when "101110000010" => data <= sine_rom(2946);
     when "101110000011" => data <= sine_rom(2947);
     when "101110000100" => data <= sine_rom(2948);
     when "101110000101" => data <= sine_rom(2949);
     when "101110000110" => data <= sine_rom(2950);
     when "101110000111" => data <= sine_rom(2951);
     when "101110001000" => data <= sine_rom(2952);
     when "101110001001" => data <= sine_rom(2953);
     when "101110001010" => data <= sine_rom(2954);
     when "101110001011" => data <= sine_rom(2955);
     when "101110001100" => data <= sine_rom(2956);
     when "101110001101" => data <= sine_rom(2957);
     when "101110001110" => data <= sine_rom(2958);
     when "101110001111" => data <= sine_rom(2959);
     when "101110010000" => data <= sine_rom(2960);
     when "101110010001" => data <= sine_rom(2961);
     when "101110010010" => data <= sine_rom(2962);
     when "101110010011" => data <= sine_rom(2963);
     when "101110010100" => data <= sine_rom(2964);
     when "101110010101" => data <= sine_rom(2965);
     when "101110010110" => data <= sine_rom(2966);
     when "101110010111" => data <= sine_rom(2967);
     when "101110011000" => data <= sine_rom(2968);
     when "101110011001" => data <= sine_rom(2969);
     when "101110011010" => data <= sine_rom(2970);
     when "101110011011" => data <= sine_rom(2971);
     when "101110011100" => data <= sine_rom(2972);
     when "101110011101" => data <= sine_rom(2973);
     when "101110011110" => data <= sine_rom(2974);
     when "101110011111" => data <= sine_rom(2975);
     when "101110100000" => data <= sine_rom(2976);
     when "101110100001" => data <= sine_rom(2977);
     when "101110100010" => data <= sine_rom(2978);
     when "101110100011" => data <= sine_rom(2979);
     when "101110100100" => data <= sine_rom(2980);
     when "101110100101" => data <= sine_rom(2981);
     when "101110100110" => data <= sine_rom(2982);
     when "101110100111" => data <= sine_rom(2983);
     when "101110101000" => data <= sine_rom(2984);
     when "101110101001" => data <= sine_rom(2985);
     when "101110101010" => data <= sine_rom(2986);
     when "101110101011" => data <= sine_rom(2987);
     when "101110101100" => data <= sine_rom(2988);
     when "101110101101" => data <= sine_rom(2989);
     when "101110101110" => data <= sine_rom(2990);
     when "101110101111" => data <= sine_rom(2991);
     when "101110110000" => data <= sine_rom(2992);
     when "101110110001" => data <= sine_rom(2993);
     when "101110110010" => data <= sine_rom(2994);
     when "101110110011" => data <= sine_rom(2995);
     when "101110110100" => data <= sine_rom(2996);
     when "101110110101" => data <= sine_rom(2997);
     when "101110110110" => data <= sine_rom(2998);
     when "101110110111" => data <= sine_rom(2999);
     when "101110111000" => data <= sine_rom(3000);
     when "101110111001" => data <= sine_rom(3001);
     when "101110111010" => data <= sine_rom(3002);
     when "101110111011" => data <= sine_rom(3003);
     when "101110111100" => data <= sine_rom(3004);
     when "101110111101" => data <= sine_rom(3005);
     when "101110111110" => data <= sine_rom(3006);
     when "101110111111" => data <= sine_rom(3007);
     when "101111000000" => data <= sine_rom(3008);
     when "101111000001" => data <= sine_rom(3009);
     when "101111000010" => data <= sine_rom(3010);
     when "101111000011" => data <= sine_rom(3011);
     when "101111000100" => data <= sine_rom(3012);
     when "101111000101" => data <= sine_rom(3013);
     when "101111000110" => data <= sine_rom(3014);
     when "101111000111" => data <= sine_rom(3015);
     when "101111001000" => data <= sine_rom(3016);
     when "101111001001" => data <= sine_rom(3017);
     when "101111001010" => data <= sine_rom(3018);
     when "101111001011" => data <= sine_rom(3019);
     when "101111001100" => data <= sine_rom(3020);
     when "101111001101" => data <= sine_rom(3021);
     when "101111001110" => data <= sine_rom(3022);
     when "101111001111" => data <= sine_rom(3023);
     when "101111010000" => data <= sine_rom(3024);
     when "101111010001" => data <= sine_rom(3025);
     when "101111010010" => data <= sine_rom(3026);
     when "101111010011" => data <= sine_rom(3027);
     when "101111010100" => data <= sine_rom(3028);
     when "101111010101" => data <= sine_rom(3029);
     when "101111010110" => data <= sine_rom(3030);
     when "101111010111" => data <= sine_rom(3031);
     when "101111011000" => data <= sine_rom(3032);
     when "101111011001" => data <= sine_rom(3033);
     when "101111011010" => data <= sine_rom(3034);
     when "101111011011" => data <= sine_rom(3035);
     when "101111011100" => data <= sine_rom(3036);
     when "101111011101" => data <= sine_rom(3037);
     when "101111011110" => data <= sine_rom(3038);
     when "101111011111" => data <= sine_rom(3039);
     when "101111100000" => data <= sine_rom(3040);
     when "101111100001" => data <= sine_rom(3041);
     when "101111100010" => data <= sine_rom(3042);
     when "101111100011" => data <= sine_rom(3043);
     when "101111100100" => data <= sine_rom(3044);
     when "101111100101" => data <= sine_rom(3045);
     when "101111100110" => data <= sine_rom(3046);
     when "101111100111" => data <= sine_rom(3047);
     when "101111101000" => data <= sine_rom(3048);
     when "101111101001" => data <= sine_rom(3049);
     when "101111101010" => data <= sine_rom(3050);
     when "101111101011" => data <= sine_rom(3051);
     when "101111101100" => data <= sine_rom(3052);
     when "101111101101" => data <= sine_rom(3053);
     when "101111101110" => data <= sine_rom(3054);
     when "101111101111" => data <= sine_rom(3055);
     when "101111110000" => data <= sine_rom(3056);
     when "101111110001" => data <= sine_rom(3057);
     when "101111110010" => data <= sine_rom(3058);
     when "101111110011" => data <= sine_rom(3059);
     when "101111110100" => data <= sine_rom(3060);
     when "101111110101" => data <= sine_rom(3061);
     when "101111110110" => data <= sine_rom(3062);
     when "101111110111" => data <= sine_rom(3063);
     when "101111111000" => data <= sine_rom(3064);
     when "101111111001" => data <= sine_rom(3065);
     when "101111111010" => data <= sine_rom(3066);
     when "101111111011" => data <= sine_rom(3067);
     when "101111111100" => data <= sine_rom(3068);
     when "101111111101" => data <= sine_rom(3069);
     when "101111111110" => data <= sine_rom(3070);
     when "101111111111" => data <= sine_rom(3071);
     when "110000000000" => data <= sine_rom(3072);
     when "110000000001" => data <= sine_rom(3073);
     when "110000000010" => data <= sine_rom(3074);
     when "110000000011" => data <= sine_rom(3075);
     when "110000000100" => data <= sine_rom(3076);
     when "110000000101" => data <= sine_rom(3077);
     when "110000000110" => data <= sine_rom(3078);
     when "110000000111" => data <= sine_rom(3079);
     when "110000001000" => data <= sine_rom(3080);
     when "110000001001" => data <= sine_rom(3081);
     when "110000001010" => data <= sine_rom(3082);
     when "110000001011" => data <= sine_rom(3083);
     when "110000001100" => data <= sine_rom(3084);
     when "110000001101" => data <= sine_rom(3085);
     when "110000001110" => data <= sine_rom(3086);
     when "110000001111" => data <= sine_rom(3087);
     when "110000010000" => data <= sine_rom(3088);
     when "110000010001" => data <= sine_rom(3089);
     when "110000010010" => data <= sine_rom(3090);
     when "110000010011" => data <= sine_rom(3091);
     when "110000010100" => data <= sine_rom(3092);
     when "110000010101" => data <= sine_rom(3093);
     when "110000010110" => data <= sine_rom(3094);
     when "110000010111" => data <= sine_rom(3095);
     when "110000011000" => data <= sine_rom(3096);
     when "110000011001" => data <= sine_rom(3097);
     when "110000011010" => data <= sine_rom(3098);
     when "110000011011" => data <= sine_rom(3099);
     when "110000011100" => data <= sine_rom(3100);
     when "110000011101" => data <= sine_rom(3101);
     when "110000011110" => data <= sine_rom(3102);
     when "110000011111" => data <= sine_rom(3103);
     when "110000100000" => data <= sine_rom(3104);
     when "110000100001" => data <= sine_rom(3105);
     when "110000100010" => data <= sine_rom(3106);
     when "110000100011" => data <= sine_rom(3107);
     when "110000100100" => data <= sine_rom(3108);
     when "110000100101" => data <= sine_rom(3109);
     when "110000100110" => data <= sine_rom(3110);
     when "110000100111" => data <= sine_rom(3111);
     when "110000101000" => data <= sine_rom(3112);
     when "110000101001" => data <= sine_rom(3113);
     when "110000101010" => data <= sine_rom(3114);
     when "110000101011" => data <= sine_rom(3115);
     when "110000101100" => data <= sine_rom(3116);
     when "110000101101" => data <= sine_rom(3117);
     when "110000101110" => data <= sine_rom(3118);
     when "110000101111" => data <= sine_rom(3119);
     when "110000110000" => data <= sine_rom(3120);
     when "110000110001" => data <= sine_rom(3121);
     when "110000110010" => data <= sine_rom(3122);
     when "110000110011" => data <= sine_rom(3123);
     when "110000110100" => data <= sine_rom(3124);
     when "110000110101" => data <= sine_rom(3125);
     when "110000110110" => data <= sine_rom(3126);
     when "110000110111" => data <= sine_rom(3127);
     when "110000111000" => data <= sine_rom(3128);
     when "110000111001" => data <= sine_rom(3129);
     when "110000111010" => data <= sine_rom(3130);
     when "110000111011" => data <= sine_rom(3131);
     when "110000111100" => data <= sine_rom(3132);
     when "110000111101" => data <= sine_rom(3133);
     when "110000111110" => data <= sine_rom(3134);
     when "110000111111" => data <= sine_rom(3135);
     when "110001000000" => data <= sine_rom(3136);
     when "110001000001" => data <= sine_rom(3137);
     when "110001000010" => data <= sine_rom(3138);
     when "110001000011" => data <= sine_rom(3139);
     when "110001000100" => data <= sine_rom(3140);
     when "110001000101" => data <= sine_rom(3141);
     when "110001000110" => data <= sine_rom(3142);
     when "110001000111" => data <= sine_rom(3143);
     when "110001001000" => data <= sine_rom(3144);
     when "110001001001" => data <= sine_rom(3145);
     when "110001001010" => data <= sine_rom(3146);
     when "110001001011" => data <= sine_rom(3147);
     when "110001001100" => data <= sine_rom(3148);
     when "110001001101" => data <= sine_rom(3149);
     when "110001001110" => data <= sine_rom(3150);
     when "110001001111" => data <= sine_rom(3151);
     when "110001010000" => data <= sine_rom(3152);
     when "110001010001" => data <= sine_rom(3153);
     when "110001010010" => data <= sine_rom(3154);
     when "110001010011" => data <= sine_rom(3155);
     when "110001010100" => data <= sine_rom(3156);
     when "110001010101" => data <= sine_rom(3157);
     when "110001010110" => data <= sine_rom(3158);
     when "110001010111" => data <= sine_rom(3159);
     when "110001011000" => data <= sine_rom(3160);
     when "110001011001" => data <= sine_rom(3161);
     when "110001011010" => data <= sine_rom(3162);
     when "110001011011" => data <= sine_rom(3163);
     when "110001011100" => data <= sine_rom(3164);
     when "110001011101" => data <= sine_rom(3165);
     when "110001011110" => data <= sine_rom(3166);
     when "110001011111" => data <= sine_rom(3167);
     when "110001100000" => data <= sine_rom(3168);
     when "110001100001" => data <= sine_rom(3169);
     when "110001100010" => data <= sine_rom(3170);
     when "110001100011" => data <= sine_rom(3171);
     when "110001100100" => data <= sine_rom(3172);
     when "110001100101" => data <= sine_rom(3173);
     when "110001100110" => data <= sine_rom(3174);
     when "110001100111" => data <= sine_rom(3175);
     when "110001101000" => data <= sine_rom(3176);
     when "110001101001" => data <= sine_rom(3177);
     when "110001101010" => data <= sine_rom(3178);
     when "110001101011" => data <= sine_rom(3179);
     when "110001101100" => data <= sine_rom(3180);
     when "110001101101" => data <= sine_rom(3181);
     when "110001101110" => data <= sine_rom(3182);
     when "110001101111" => data <= sine_rom(3183);
     when "110001110000" => data <= sine_rom(3184);
     when "110001110001" => data <= sine_rom(3185);
     when "110001110010" => data <= sine_rom(3186);
     when "110001110011" => data <= sine_rom(3187);
     when "110001110100" => data <= sine_rom(3188);
     when "110001110101" => data <= sine_rom(3189);
     when "110001110110" => data <= sine_rom(3190);
     when "110001110111" => data <= sine_rom(3191);
     when "110001111000" => data <= sine_rom(3192);
     when "110001111001" => data <= sine_rom(3193);
     when "110001111010" => data <= sine_rom(3194);
     when "110001111011" => data <= sine_rom(3195);
     when "110001111100" => data <= sine_rom(3196);
     when "110001111101" => data <= sine_rom(3197);
     when "110001111110" => data <= sine_rom(3198);
     when "110001111111" => data <= sine_rom(3199);
     when "110010000000" => data <= sine_rom(3200);
     when "110010000001" => data <= sine_rom(3201);
     when "110010000010" => data <= sine_rom(3202);
     when "110010000011" => data <= sine_rom(3203);
     when "110010000100" => data <= sine_rom(3204);
     when "110010000101" => data <= sine_rom(3205);
     when "110010000110" => data <= sine_rom(3206);
     when "110010000111" => data <= sine_rom(3207);
     when "110010001000" => data <= sine_rom(3208);
     when "110010001001" => data <= sine_rom(3209);
     when "110010001010" => data <= sine_rom(3210);
     when "110010001011" => data <= sine_rom(3211);
     when "110010001100" => data <= sine_rom(3212);
     when "110010001101" => data <= sine_rom(3213);
     when "110010001110" => data <= sine_rom(3214);
     when "110010001111" => data <= sine_rom(3215);
     when "110010010000" => data <= sine_rom(3216);
     when "110010010001" => data <= sine_rom(3217);
     when "110010010010" => data <= sine_rom(3218);
     when "110010010011" => data <= sine_rom(3219);
     when "110010010100" => data <= sine_rom(3220);
     when "110010010101" => data <= sine_rom(3221);
     when "110010010110" => data <= sine_rom(3222);
     when "110010010111" => data <= sine_rom(3223);
     when "110010011000" => data <= sine_rom(3224);
     when "110010011001" => data <= sine_rom(3225);
     when "110010011010" => data <= sine_rom(3226);
     when "110010011011" => data <= sine_rom(3227);
     when "110010011100" => data <= sine_rom(3228);
     when "110010011101" => data <= sine_rom(3229);
     when "110010011110" => data <= sine_rom(3230);
     when "110010011111" => data <= sine_rom(3231);
     when "110010100000" => data <= sine_rom(3232);
     when "110010100001" => data <= sine_rom(3233);
     when "110010100010" => data <= sine_rom(3234);
     when "110010100011" => data <= sine_rom(3235);
     when "110010100100" => data <= sine_rom(3236);
     when "110010100101" => data <= sine_rom(3237);
     when "110010100110" => data <= sine_rom(3238);
     when "110010100111" => data <= sine_rom(3239);
     when "110010101000" => data <= sine_rom(3240);
     when "110010101001" => data <= sine_rom(3241);
     when "110010101010" => data <= sine_rom(3242);
     when "110010101011" => data <= sine_rom(3243);
     when "110010101100" => data <= sine_rom(3244);
     when "110010101101" => data <= sine_rom(3245);
     when "110010101110" => data <= sine_rom(3246);
     when "110010101111" => data <= sine_rom(3247);
     when "110010110000" => data <= sine_rom(3248);
     when "110010110001" => data <= sine_rom(3249);
     when "110010110010" => data <= sine_rom(3250);
     when "110010110011" => data <= sine_rom(3251);
     when "110010110100" => data <= sine_rom(3252);
     when "110010110101" => data <= sine_rom(3253);
     when "110010110110" => data <= sine_rom(3254);
     when "110010110111" => data <= sine_rom(3255);
     when "110010111000" => data <= sine_rom(3256);
     when "110010111001" => data <= sine_rom(3257);
     when "110010111010" => data <= sine_rom(3258);
     when "110010111011" => data <= sine_rom(3259);
     when "110010111100" => data <= sine_rom(3260);
     when "110010111101" => data <= sine_rom(3261);
     when "110010111110" => data <= sine_rom(3262);
     when "110010111111" => data <= sine_rom(3263);
     when "110011000000" => data <= sine_rom(3264);
     when "110011000001" => data <= sine_rom(3265);
     when "110011000010" => data <= sine_rom(3266);
     when "110011000011" => data <= sine_rom(3267);
     when "110011000100" => data <= sine_rom(3268);
     when "110011000101" => data <= sine_rom(3269);
     when "110011000110" => data <= sine_rom(3270);
     when "110011000111" => data <= sine_rom(3271);
     when "110011001000" => data <= sine_rom(3272);
     when "110011001001" => data <= sine_rom(3273);
     when "110011001010" => data <= sine_rom(3274);
     when "110011001011" => data <= sine_rom(3275);
     when "110011001100" => data <= sine_rom(3276);
     when "110011001101" => data <= sine_rom(3277);
     when "110011001110" => data <= sine_rom(3278);
     when "110011001111" => data <= sine_rom(3279);
     when "110011010000" => data <= sine_rom(3280);
     when "110011010001" => data <= sine_rom(3281);
     when "110011010010" => data <= sine_rom(3282);
     when "110011010011" => data <= sine_rom(3283);
     when "110011010100" => data <= sine_rom(3284);
     when "110011010101" => data <= sine_rom(3285);
     when "110011010110" => data <= sine_rom(3286);
     when "110011010111" => data <= sine_rom(3287);
     when "110011011000" => data <= sine_rom(3288);
     when "110011011001" => data <= sine_rom(3289);
     when "110011011010" => data <= sine_rom(3290);
     when "110011011011" => data <= sine_rom(3291);
     when "110011011100" => data <= sine_rom(3292);
     when "110011011101" => data <= sine_rom(3293);
     when "110011011110" => data <= sine_rom(3294);
     when "110011011111" => data <= sine_rom(3295);
     when "110011100000" => data <= sine_rom(3296);
     when "110011100001" => data <= sine_rom(3297);
     when "110011100010" => data <= sine_rom(3298);
     when "110011100011" => data <= sine_rom(3299);
     when "110011100100" => data <= sine_rom(3300);
     when "110011100101" => data <= sine_rom(3301);
     when "110011100110" => data <= sine_rom(3302);
     when "110011100111" => data <= sine_rom(3303);
     when "110011101000" => data <= sine_rom(3304);
     when "110011101001" => data <= sine_rom(3305);
     when "110011101010" => data <= sine_rom(3306);
     when "110011101011" => data <= sine_rom(3307);
     when "110011101100" => data <= sine_rom(3308);
     when "110011101101" => data <= sine_rom(3309);
     when "110011101110" => data <= sine_rom(3310);
     when "110011101111" => data <= sine_rom(3311);
     when "110011110000" => data <= sine_rom(3312);
     when "110011110001" => data <= sine_rom(3313);
     when "110011110010" => data <= sine_rom(3314);
     when "110011110011" => data <= sine_rom(3315);
     when "110011110100" => data <= sine_rom(3316);
     when "110011110101" => data <= sine_rom(3317);
     when "110011110110" => data <= sine_rom(3318);
     when "110011110111" => data <= sine_rom(3319);
     when "110011111000" => data <= sine_rom(3320);
     when "110011111001" => data <= sine_rom(3321);
     when "110011111010" => data <= sine_rom(3322);
     when "110011111011" => data <= sine_rom(3323);
     when "110011111100" => data <= sine_rom(3324);
     when "110011111101" => data <= sine_rom(3325);
     when "110011111110" => data <= sine_rom(3326);
     when "110011111111" => data <= sine_rom(3327);
     when "110100000000" => data <= sine_rom(3328);
     when "110100000001" => data <= sine_rom(3329);
     when "110100000010" => data <= sine_rom(3330);
     when "110100000011" => data <= sine_rom(3331);
     when "110100000100" => data <= sine_rom(3332);
     when "110100000101" => data <= sine_rom(3333);
     when "110100000110" => data <= sine_rom(3334);
     when "110100000111" => data <= sine_rom(3335);
     when "110100001000" => data <= sine_rom(3336);
     when "110100001001" => data <= sine_rom(3337);
     when "110100001010" => data <= sine_rom(3338);
     when "110100001011" => data <= sine_rom(3339);
     when "110100001100" => data <= sine_rom(3340);
     when "110100001101" => data <= sine_rom(3341);
     when "110100001110" => data <= sine_rom(3342);
     when "110100001111" => data <= sine_rom(3343);
     when "110100010000" => data <= sine_rom(3344);
     when "110100010001" => data <= sine_rom(3345);
     when "110100010010" => data <= sine_rom(3346);
     when "110100010011" => data <= sine_rom(3347);
     when "110100010100" => data <= sine_rom(3348);
     when "110100010101" => data <= sine_rom(3349);
     when "110100010110" => data <= sine_rom(3350);
     when "110100010111" => data <= sine_rom(3351);
     when "110100011000" => data <= sine_rom(3352);
     when "110100011001" => data <= sine_rom(3353);
     when "110100011010" => data <= sine_rom(3354);
     when "110100011011" => data <= sine_rom(3355);
     when "110100011100" => data <= sine_rom(3356);
     when "110100011101" => data <= sine_rom(3357);
     when "110100011110" => data <= sine_rom(3358);
     when "110100011111" => data <= sine_rom(3359);
     when "110100100000" => data <= sine_rom(3360);
     when "110100100001" => data <= sine_rom(3361);
     when "110100100010" => data <= sine_rom(3362);
     when "110100100011" => data <= sine_rom(3363);
     when "110100100100" => data <= sine_rom(3364);
     when "110100100101" => data <= sine_rom(3365);
     when "110100100110" => data <= sine_rom(3366);
     when "110100100111" => data <= sine_rom(3367);
     when "110100101000" => data <= sine_rom(3368);
     when "110100101001" => data <= sine_rom(3369);
     when "110100101010" => data <= sine_rom(3370);
     when "110100101011" => data <= sine_rom(3371);
     when "110100101100" => data <= sine_rom(3372);
     when "110100101101" => data <= sine_rom(3373);
     when "110100101110" => data <= sine_rom(3374);
     when "110100101111" => data <= sine_rom(3375);
     when "110100110000" => data <= sine_rom(3376);
     when "110100110001" => data <= sine_rom(3377);
     when "110100110010" => data <= sine_rom(3378);
     when "110100110011" => data <= sine_rom(3379);
     when "110100110100" => data <= sine_rom(3380);
     when "110100110101" => data <= sine_rom(3381);
     when "110100110110" => data <= sine_rom(3382);
     when "110100110111" => data <= sine_rom(3383);
     when "110100111000" => data <= sine_rom(3384);
     when "110100111001" => data <= sine_rom(3385);
     when "110100111010" => data <= sine_rom(3386);
     when "110100111011" => data <= sine_rom(3387);
     when "110100111100" => data <= sine_rom(3388);
     when "110100111101" => data <= sine_rom(3389);
     when "110100111110" => data <= sine_rom(3390);
     when "110100111111" => data <= sine_rom(3391);
     when "110101000000" => data <= sine_rom(3392);
     when "110101000001" => data <= sine_rom(3393);
     when "110101000010" => data <= sine_rom(3394);
     when "110101000011" => data <= sine_rom(3395);
     when "110101000100" => data <= sine_rom(3396);
     when "110101000101" => data <= sine_rom(3397);
     when "110101000110" => data <= sine_rom(3398);
     when "110101000111" => data <= sine_rom(3399);
     when "110101001000" => data <= sine_rom(3400);
     when "110101001001" => data <= sine_rom(3401);
     when "110101001010" => data <= sine_rom(3402);
     when "110101001011" => data <= sine_rom(3403);
     when "110101001100" => data <= sine_rom(3404);
     when "110101001101" => data <= sine_rom(3405);
     when "110101001110" => data <= sine_rom(3406);
     when "110101001111" => data <= sine_rom(3407);
     when "110101010000" => data <= sine_rom(3408);
     when "110101010001" => data <= sine_rom(3409);
     when "110101010010" => data <= sine_rom(3410);
     when "110101010011" => data <= sine_rom(3411);
     when "110101010100" => data <= sine_rom(3412);
     when "110101010101" => data <= sine_rom(3413);
     when "110101010110" => data <= sine_rom(3414);
     when "110101010111" => data <= sine_rom(3415);
     when "110101011000" => data <= sine_rom(3416);
     when "110101011001" => data <= sine_rom(3417);
     when "110101011010" => data <= sine_rom(3418);
     when "110101011011" => data <= sine_rom(3419);
     when "110101011100" => data <= sine_rom(3420);
     when "110101011101" => data <= sine_rom(3421);
     when "110101011110" => data <= sine_rom(3422);
     when "110101011111" => data <= sine_rom(3423);
     when "110101100000" => data <= sine_rom(3424);
     when "110101100001" => data <= sine_rom(3425);
     when "110101100010" => data <= sine_rom(3426);
     when "110101100011" => data <= sine_rom(3427);
     when "110101100100" => data <= sine_rom(3428);
     when "110101100101" => data <= sine_rom(3429);
     when "110101100110" => data <= sine_rom(3430);
     when "110101100111" => data <= sine_rom(3431);
     when "110101101000" => data <= sine_rom(3432);
     when "110101101001" => data <= sine_rom(3433);
     when "110101101010" => data <= sine_rom(3434);
     when "110101101011" => data <= sine_rom(3435);
     when "110101101100" => data <= sine_rom(3436);
     when "110101101101" => data <= sine_rom(3437);
     when "110101101110" => data <= sine_rom(3438);
     when "110101101111" => data <= sine_rom(3439);
     when "110101110000" => data <= sine_rom(3440);
     when "110101110001" => data <= sine_rom(3441);
     when "110101110010" => data <= sine_rom(3442);
     when "110101110011" => data <= sine_rom(3443);
     when "110101110100" => data <= sine_rom(3444);
     when "110101110101" => data <= sine_rom(3445);
     when "110101110110" => data <= sine_rom(3446);
     when "110101110111" => data <= sine_rom(3447);
     when "110101111000" => data <= sine_rom(3448);
     when "110101111001" => data <= sine_rom(3449);
     when "110101111010" => data <= sine_rom(3450);
     when "110101111011" => data <= sine_rom(3451);
     when "110101111100" => data <= sine_rom(3452);
     when "110101111101" => data <= sine_rom(3453);
     when "110101111110" => data <= sine_rom(3454);
     when "110101111111" => data <= sine_rom(3455);
     when "110110000000" => data <= sine_rom(3456);
     when "110110000001" => data <= sine_rom(3457);
     when "110110000010" => data <= sine_rom(3458);
     when "110110000011" => data <= sine_rom(3459);
     when "110110000100" => data <= sine_rom(3460);
     when "110110000101" => data <= sine_rom(3461);
     when "110110000110" => data <= sine_rom(3462);
     when "110110000111" => data <= sine_rom(3463);
     when "110110001000" => data <= sine_rom(3464);
     when "110110001001" => data <= sine_rom(3465);
     when "110110001010" => data <= sine_rom(3466);
     when "110110001011" => data <= sine_rom(3467);
     when "110110001100" => data <= sine_rom(3468);
     when "110110001101" => data <= sine_rom(3469);
     when "110110001110" => data <= sine_rom(3470);
     when "110110001111" => data <= sine_rom(3471);
     when "110110010000" => data <= sine_rom(3472);
     when "110110010001" => data <= sine_rom(3473);
     when "110110010010" => data <= sine_rom(3474);
     when "110110010011" => data <= sine_rom(3475);
     when "110110010100" => data <= sine_rom(3476);
     when "110110010101" => data <= sine_rom(3477);
     when "110110010110" => data <= sine_rom(3478);
     when "110110010111" => data <= sine_rom(3479);
     when "110110011000" => data <= sine_rom(3480);
     when "110110011001" => data <= sine_rom(3481);
     when "110110011010" => data <= sine_rom(3482);
     when "110110011011" => data <= sine_rom(3483);
     when "110110011100" => data <= sine_rom(3484);
     when "110110011101" => data <= sine_rom(3485);
     when "110110011110" => data <= sine_rom(3486);
     when "110110011111" => data <= sine_rom(3487);
     when "110110100000" => data <= sine_rom(3488);
     when "110110100001" => data <= sine_rom(3489);
     when "110110100010" => data <= sine_rom(3490);
     when "110110100011" => data <= sine_rom(3491);
     when "110110100100" => data <= sine_rom(3492);
     when "110110100101" => data <= sine_rom(3493);
     when "110110100110" => data <= sine_rom(3494);
     when "110110100111" => data <= sine_rom(3495);
     when "110110101000" => data <= sine_rom(3496);
     when "110110101001" => data <= sine_rom(3497);
     when "110110101010" => data <= sine_rom(3498);
     when "110110101011" => data <= sine_rom(3499);
     when "110110101100" => data <= sine_rom(3500);
     when "110110101101" => data <= sine_rom(3501);
     when "110110101110" => data <= sine_rom(3502);
     when "110110101111" => data <= sine_rom(3503);
     when "110110110000" => data <= sine_rom(3504);
     when "110110110001" => data <= sine_rom(3505);
     when "110110110010" => data <= sine_rom(3506);
     when "110110110011" => data <= sine_rom(3507);
     when "110110110100" => data <= sine_rom(3508);
     when "110110110101" => data <= sine_rom(3509);
     when "110110110110" => data <= sine_rom(3510);
     when "110110110111" => data <= sine_rom(3511);
     when "110110111000" => data <= sine_rom(3512);
     when "110110111001" => data <= sine_rom(3513);
     when "110110111010" => data <= sine_rom(3514);
     when "110110111011" => data <= sine_rom(3515);
     when "110110111100" => data <= sine_rom(3516);
     when "110110111101" => data <= sine_rom(3517);
     when "110110111110" => data <= sine_rom(3518);
     when "110110111111" => data <= sine_rom(3519);
     when "110111000000" => data <= sine_rom(3520);
     when "110111000001" => data <= sine_rom(3521);
     when "110111000010" => data <= sine_rom(3522);
     when "110111000011" => data <= sine_rom(3523);
     when "110111000100" => data <= sine_rom(3524);
     when "110111000101" => data <= sine_rom(3525);
     when "110111000110" => data <= sine_rom(3526);
     when "110111000111" => data <= sine_rom(3527);
     when "110111001000" => data <= sine_rom(3528);
     when "110111001001" => data <= sine_rom(3529);
     when "110111001010" => data <= sine_rom(3530);
     when "110111001011" => data <= sine_rom(3531);
     when "110111001100" => data <= sine_rom(3532);
     when "110111001101" => data <= sine_rom(3533);
     when "110111001110" => data <= sine_rom(3534);
     when "110111001111" => data <= sine_rom(3535);
     when "110111010000" => data <= sine_rom(3536);
     when "110111010001" => data <= sine_rom(3537);
     when "110111010010" => data <= sine_rom(3538);
     when "110111010011" => data <= sine_rom(3539);
     when "110111010100" => data <= sine_rom(3540);
     when "110111010101" => data <= sine_rom(3541);
     when "110111010110" => data <= sine_rom(3542);
     when "110111010111" => data <= sine_rom(3543);
     when "110111011000" => data <= sine_rom(3544);
     when "110111011001" => data <= sine_rom(3545);
     when "110111011010" => data <= sine_rom(3546);
     when "110111011011" => data <= sine_rom(3547);
     when "110111011100" => data <= sine_rom(3548);
     when "110111011101" => data <= sine_rom(3549);
     when "110111011110" => data <= sine_rom(3550);
     when "110111011111" => data <= sine_rom(3551);
     when "110111100000" => data <= sine_rom(3552);
     when "110111100001" => data <= sine_rom(3553);
     when "110111100010" => data <= sine_rom(3554);
     when "110111100011" => data <= sine_rom(3555);
     when "110111100100" => data <= sine_rom(3556);
     when "110111100101" => data <= sine_rom(3557);
     when "110111100110" => data <= sine_rom(3558);
     when "110111100111" => data <= sine_rom(3559);
     when "110111101000" => data <= sine_rom(3560);
     when "110111101001" => data <= sine_rom(3561);
     when "110111101010" => data <= sine_rom(3562);
     when "110111101011" => data <= sine_rom(3563);
     when "110111101100" => data <= sine_rom(3564);
     when "110111101101" => data <= sine_rom(3565);
     when "110111101110" => data <= sine_rom(3566);
     when "110111101111" => data <= sine_rom(3567);
     when "110111110000" => data <= sine_rom(3568);
     when "110111110001" => data <= sine_rom(3569);
     when "110111110010" => data <= sine_rom(3570);
     when "110111110011" => data <= sine_rom(3571);
     when "110111110100" => data <= sine_rom(3572);
     when "110111110101" => data <= sine_rom(3573);
     when "110111110110" => data <= sine_rom(3574);
     when "110111110111" => data <= sine_rom(3575);
     when "110111111000" => data <= sine_rom(3576);
     when "110111111001" => data <= sine_rom(3577);
     when "110111111010" => data <= sine_rom(3578);
     when "110111111011" => data <= sine_rom(3579);
     when "110111111100" => data <= sine_rom(3580);
     when "110111111101" => data <= sine_rom(3581);
     when "110111111110" => data <= sine_rom(3582);
     when "110111111111" => data <= sine_rom(3583);
     when "111000000000" => data <= sine_rom(3584);
     when "111000000001" => data <= sine_rom(3585);
     when "111000000010" => data <= sine_rom(3586);
     when "111000000011" => data <= sine_rom(3587);
     when "111000000100" => data <= sine_rom(3588);
     when "111000000101" => data <= sine_rom(3589);
     when "111000000110" => data <= sine_rom(3590);
     when "111000000111" => data <= sine_rom(3591);
     when "111000001000" => data <= sine_rom(3592);
     when "111000001001" => data <= sine_rom(3593);
     when "111000001010" => data <= sine_rom(3594);
     when "111000001011" => data <= sine_rom(3595);
     when "111000001100" => data <= sine_rom(3596);
     when "111000001101" => data <= sine_rom(3597);
     when "111000001110" => data <= sine_rom(3598);
     when "111000001111" => data <= sine_rom(3599);
     when "111000010000" => data <= sine_rom(3600);
     when "111000010001" => data <= sine_rom(3601);
     when "111000010010" => data <= sine_rom(3602);
     when "111000010011" => data <= sine_rom(3603);
     when "111000010100" => data <= sine_rom(3604);
     when "111000010101" => data <= sine_rom(3605);
     when "111000010110" => data <= sine_rom(3606);
     when "111000010111" => data <= sine_rom(3607);
     when "111000011000" => data <= sine_rom(3608);
     when "111000011001" => data <= sine_rom(3609);
     when "111000011010" => data <= sine_rom(3610);
     when "111000011011" => data <= sine_rom(3611);
     when "111000011100" => data <= sine_rom(3612);
     when "111000011101" => data <= sine_rom(3613);
     when "111000011110" => data <= sine_rom(3614);
     when "111000011111" => data <= sine_rom(3615);
     when "111000100000" => data <= sine_rom(3616);
     when "111000100001" => data <= sine_rom(3617);
     when "111000100010" => data <= sine_rom(3618);
     when "111000100011" => data <= sine_rom(3619);
     when "111000100100" => data <= sine_rom(3620);
     when "111000100101" => data <= sine_rom(3621);
     when "111000100110" => data <= sine_rom(3622);
     when "111000100111" => data <= sine_rom(3623);
     when "111000101000" => data <= sine_rom(3624);
     when "111000101001" => data <= sine_rom(3625);
     when "111000101010" => data <= sine_rom(3626);
     when "111000101011" => data <= sine_rom(3627);
     when "111000101100" => data <= sine_rom(3628);
     when "111000101101" => data <= sine_rom(3629);
     when "111000101110" => data <= sine_rom(3630);
     when "111000101111" => data <= sine_rom(3631);
     when "111000110000" => data <= sine_rom(3632);
     when "111000110001" => data <= sine_rom(3633);
     when "111000110010" => data <= sine_rom(3634);
     when "111000110011" => data <= sine_rom(3635);
     when "111000110100" => data <= sine_rom(3636);
     when "111000110101" => data <= sine_rom(3637);
     when "111000110110" => data <= sine_rom(3638);
     when "111000110111" => data <= sine_rom(3639);
     when "111000111000" => data <= sine_rom(3640);
     when "111000111001" => data <= sine_rom(3641);
     when "111000111010" => data <= sine_rom(3642);
     when "111000111011" => data <= sine_rom(3643);
     when "111000111100" => data <= sine_rom(3644);
     when "111000111101" => data <= sine_rom(3645);
     when "111000111110" => data <= sine_rom(3646);
     when "111000111111" => data <= sine_rom(3647);
     when "111001000000" => data <= sine_rom(3648);
     when "111001000001" => data <= sine_rom(3649);
     when "111001000010" => data <= sine_rom(3650);
     when "111001000011" => data <= sine_rom(3651);
     when "111001000100" => data <= sine_rom(3652);
     when "111001000101" => data <= sine_rom(3653);
     when "111001000110" => data <= sine_rom(3654);
     when "111001000111" => data <= sine_rom(3655);
     when "111001001000" => data <= sine_rom(3656);
     when "111001001001" => data <= sine_rom(3657);
     when "111001001010" => data <= sine_rom(3658);
     when "111001001011" => data <= sine_rom(3659);
     when "111001001100" => data <= sine_rom(3660);
     when "111001001101" => data <= sine_rom(3661);
     when "111001001110" => data <= sine_rom(3662);
     when "111001001111" => data <= sine_rom(3663);
     when "111001010000" => data <= sine_rom(3664);
     when "111001010001" => data <= sine_rom(3665);
     when "111001010010" => data <= sine_rom(3666);
     when "111001010011" => data <= sine_rom(3667);
     when "111001010100" => data <= sine_rom(3668);
     when "111001010101" => data <= sine_rom(3669);
     when "111001010110" => data <= sine_rom(3670);
     when "111001010111" => data <= sine_rom(3671);
     when "111001011000" => data <= sine_rom(3672);
     when "111001011001" => data <= sine_rom(3673);
     when "111001011010" => data <= sine_rom(3674);
     when "111001011011" => data <= sine_rom(3675);
     when "111001011100" => data <= sine_rom(3676);
     when "111001011101" => data <= sine_rom(3677);
     when "111001011110" => data <= sine_rom(3678);
     when "111001011111" => data <= sine_rom(3679);
     when "111001100000" => data <= sine_rom(3680);
     when "111001100001" => data <= sine_rom(3681);
     when "111001100010" => data <= sine_rom(3682);
     when "111001100011" => data <= sine_rom(3683);
     when "111001100100" => data <= sine_rom(3684);
     when "111001100101" => data <= sine_rom(3685);
     when "111001100110" => data <= sine_rom(3686);
     when "111001100111" => data <= sine_rom(3687);
     when "111001101000" => data <= sine_rom(3688);
     when "111001101001" => data <= sine_rom(3689);
     when "111001101010" => data <= sine_rom(3690);
     when "111001101011" => data <= sine_rom(3691);
     when "111001101100" => data <= sine_rom(3692);
     when "111001101101" => data <= sine_rom(3693);
     when "111001101110" => data <= sine_rom(3694);
     when "111001101111" => data <= sine_rom(3695);
     when "111001110000" => data <= sine_rom(3696);
     when "111001110001" => data <= sine_rom(3697);
     when "111001110010" => data <= sine_rom(3698);
     when "111001110011" => data <= sine_rom(3699);
     when "111001110100" => data <= sine_rom(3700);
     when "111001110101" => data <= sine_rom(3701);
     when "111001110110" => data <= sine_rom(3702);
     when "111001110111" => data <= sine_rom(3703);
     when "111001111000" => data <= sine_rom(3704);
     when "111001111001" => data <= sine_rom(3705);
     when "111001111010" => data <= sine_rom(3706);
     when "111001111011" => data <= sine_rom(3707);
     when "111001111100" => data <= sine_rom(3708);
     when "111001111101" => data <= sine_rom(3709);
     when "111001111110" => data <= sine_rom(3710);
     when "111001111111" => data <= sine_rom(3711);
     when "111010000000" => data <= sine_rom(3712);
     when "111010000001" => data <= sine_rom(3713);
     when "111010000010" => data <= sine_rom(3714);
     when "111010000011" => data <= sine_rom(3715);
     when "111010000100" => data <= sine_rom(3716);
     when "111010000101" => data <= sine_rom(3717);
     when "111010000110" => data <= sine_rom(3718);
     when "111010000111" => data <= sine_rom(3719);
     when "111010001000" => data <= sine_rom(3720);
     when "111010001001" => data <= sine_rom(3721);
     when "111010001010" => data <= sine_rom(3722);
     when "111010001011" => data <= sine_rom(3723);
     when "111010001100" => data <= sine_rom(3724);
     when "111010001101" => data <= sine_rom(3725);
     when "111010001110" => data <= sine_rom(3726);
     when "111010001111" => data <= sine_rom(3727);
     when "111010010000" => data <= sine_rom(3728);
     when "111010010001" => data <= sine_rom(3729);
     when "111010010010" => data <= sine_rom(3730);
     when "111010010011" => data <= sine_rom(3731);
     when "111010010100" => data <= sine_rom(3732);
     when "111010010101" => data <= sine_rom(3733);
     when "111010010110" => data <= sine_rom(3734);
     when "111010010111" => data <= sine_rom(3735);
     when "111010011000" => data <= sine_rom(3736);
     when "111010011001" => data <= sine_rom(3737);
     when "111010011010" => data <= sine_rom(3738);
     when "111010011011" => data <= sine_rom(3739);
     when "111010011100" => data <= sine_rom(3740);
     when "111010011101" => data <= sine_rom(3741);
     when "111010011110" => data <= sine_rom(3742);
     when "111010011111" => data <= sine_rom(3743);
     when "111010100000" => data <= sine_rom(3744);
     when "111010100001" => data <= sine_rom(3745);
     when "111010100010" => data <= sine_rom(3746);
     when "111010100011" => data <= sine_rom(3747);
     when "111010100100" => data <= sine_rom(3748);
     when "111010100101" => data <= sine_rom(3749);
     when "111010100110" => data <= sine_rom(3750);
     when "111010100111" => data <= sine_rom(3751);
     when "111010101000" => data <= sine_rom(3752);
     when "111010101001" => data <= sine_rom(3753);
     when "111010101010" => data <= sine_rom(3754);
     when "111010101011" => data <= sine_rom(3755);
     when "111010101100" => data <= sine_rom(3756);
     when "111010101101" => data <= sine_rom(3757);
     when "111010101110" => data <= sine_rom(3758);
     when "111010101111" => data <= sine_rom(3759);
     when "111010110000" => data <= sine_rom(3760);
     when "111010110001" => data <= sine_rom(3761);
     when "111010110010" => data <= sine_rom(3762);
     when "111010110011" => data <= sine_rom(3763);
     when "111010110100" => data <= sine_rom(3764);
     when "111010110101" => data <= sine_rom(3765);
     when "111010110110" => data <= sine_rom(3766);
     when "111010110111" => data <= sine_rom(3767);
     when "111010111000" => data <= sine_rom(3768);
     when "111010111001" => data <= sine_rom(3769);
     when "111010111010" => data <= sine_rom(3770);
     when "111010111011" => data <= sine_rom(3771);
     when "111010111100" => data <= sine_rom(3772);
     when "111010111101" => data <= sine_rom(3773);
     when "111010111110" => data <= sine_rom(3774);
     when "111010111111" => data <= sine_rom(3775);
     when "111011000000" => data <= sine_rom(3776);
     when "111011000001" => data <= sine_rom(3777);
     when "111011000010" => data <= sine_rom(3778);
     when "111011000011" => data <= sine_rom(3779);
     when "111011000100" => data <= sine_rom(3780);
     when "111011000101" => data <= sine_rom(3781);
     when "111011000110" => data <= sine_rom(3782);
     when "111011000111" => data <= sine_rom(3783);
     when "111011001000" => data <= sine_rom(3784);
     when "111011001001" => data <= sine_rom(3785);
     when "111011001010" => data <= sine_rom(3786);
     when "111011001011" => data <= sine_rom(3787);
     when "111011001100" => data <= sine_rom(3788);
     when "111011001101" => data <= sine_rom(3789);
     when "111011001110" => data <= sine_rom(3790);
     when "111011001111" => data <= sine_rom(3791);
     when "111011010000" => data <= sine_rom(3792);
     when "111011010001" => data <= sine_rom(3793);
     when "111011010010" => data <= sine_rom(3794);
     when "111011010011" => data <= sine_rom(3795);
     when "111011010100" => data <= sine_rom(3796);
     when "111011010101" => data <= sine_rom(3797);
     when "111011010110" => data <= sine_rom(3798);
     when "111011010111" => data <= sine_rom(3799);
     when "111011011000" => data <= sine_rom(3800);
     when "111011011001" => data <= sine_rom(3801);
     when "111011011010" => data <= sine_rom(3802);
     when "111011011011" => data <= sine_rom(3803);
     when "111011011100" => data <= sine_rom(3804);
     when "111011011101" => data <= sine_rom(3805);
     when "111011011110" => data <= sine_rom(3806);
     when "111011011111" => data <= sine_rom(3807);
     when "111011100000" => data <= sine_rom(3808);
     when "111011100001" => data <= sine_rom(3809);
     when "111011100010" => data <= sine_rom(3810);
     when "111011100011" => data <= sine_rom(3811);
     when "111011100100" => data <= sine_rom(3812);
     when "111011100101" => data <= sine_rom(3813);
     when "111011100110" => data <= sine_rom(3814);
     when "111011100111" => data <= sine_rom(3815);
     when "111011101000" => data <= sine_rom(3816);
     when "111011101001" => data <= sine_rom(3817);
     when "111011101010" => data <= sine_rom(3818);
     when "111011101011" => data <= sine_rom(3819);
     when "111011101100" => data <= sine_rom(3820);
     when "111011101101" => data <= sine_rom(3821);
     when "111011101110" => data <= sine_rom(3822);
     when "111011101111" => data <= sine_rom(3823);
     when "111011110000" => data <= sine_rom(3824);
     when "111011110001" => data <= sine_rom(3825);
     when "111011110010" => data <= sine_rom(3826);
     when "111011110011" => data <= sine_rom(3827);
     when "111011110100" => data <= sine_rom(3828);
     when "111011110101" => data <= sine_rom(3829);
     when "111011110110" => data <= sine_rom(3830);
     when "111011110111" => data <= sine_rom(3831);
     when "111011111000" => data <= sine_rom(3832);
     when "111011111001" => data <= sine_rom(3833);
     when "111011111010" => data <= sine_rom(3834);
     when "111011111011" => data <= sine_rom(3835);
     when "111011111100" => data <= sine_rom(3836);
     when "111011111101" => data <= sine_rom(3837);
     when "111011111110" => data <= sine_rom(3838);
     when "111011111111" => data <= sine_rom(3839);
     when "111100000000" => data <= sine_rom(3840);
     when "111100000001" => data <= sine_rom(3841);
     when "111100000010" => data <= sine_rom(3842);
     when "111100000011" => data <= sine_rom(3843);
     when "111100000100" => data <= sine_rom(3844);
     when "111100000101" => data <= sine_rom(3845);
     when "111100000110" => data <= sine_rom(3846);
     when "111100000111" => data <= sine_rom(3847);
     when "111100001000" => data <= sine_rom(3848);
     when "111100001001" => data <= sine_rom(3849);
     when "111100001010" => data <= sine_rom(3850);
     when "111100001011" => data <= sine_rom(3851);
     when "111100001100" => data <= sine_rom(3852);
     when "111100001101" => data <= sine_rom(3853);
     when "111100001110" => data <= sine_rom(3854);
     when "111100001111" => data <= sine_rom(3855);
     when "111100010000" => data <= sine_rom(3856);
     when "111100010001" => data <= sine_rom(3857);
     when "111100010010" => data <= sine_rom(3858);
     when "111100010011" => data <= sine_rom(3859);
     when "111100010100" => data <= sine_rom(3860);
     when "111100010101" => data <= sine_rom(3861);
     when "111100010110" => data <= sine_rom(3862);
     when "111100010111" => data <= sine_rom(3863);
     when "111100011000" => data <= sine_rom(3864);
     when "111100011001" => data <= sine_rom(3865);
     when "111100011010" => data <= sine_rom(3866);
     when "111100011011" => data <= sine_rom(3867);
     when "111100011100" => data <= sine_rom(3868);
     when "111100011101" => data <= sine_rom(3869);
     when "111100011110" => data <= sine_rom(3870);
     when "111100011111" => data <= sine_rom(3871);
     when "111100100000" => data <= sine_rom(3872);
     when "111100100001" => data <= sine_rom(3873);
     when "111100100010" => data <= sine_rom(3874);
     when "111100100011" => data <= sine_rom(3875);
     when "111100100100" => data <= sine_rom(3876);
     when "111100100101" => data <= sine_rom(3877);
     when "111100100110" => data <= sine_rom(3878);
     when "111100100111" => data <= sine_rom(3879);
     when "111100101000" => data <= sine_rom(3880);
     when "111100101001" => data <= sine_rom(3881);
     when "111100101010" => data <= sine_rom(3882);
     when "111100101011" => data <= sine_rom(3883);
     when "111100101100" => data <= sine_rom(3884);
     when "111100101101" => data <= sine_rom(3885);
     when "111100101110" => data <= sine_rom(3886);
     when "111100101111" => data <= sine_rom(3887);
     when "111100110000" => data <= sine_rom(3888);
     when "111100110001" => data <= sine_rom(3889);
     when "111100110010" => data <= sine_rom(3890);
     when "111100110011" => data <= sine_rom(3891);
     when "111100110100" => data <= sine_rom(3892);
     when "111100110101" => data <= sine_rom(3893);
     when "111100110110" => data <= sine_rom(3894);
     when "111100110111" => data <= sine_rom(3895);
     when "111100111000" => data <= sine_rom(3896);
     when "111100111001" => data <= sine_rom(3897);
     when "111100111010" => data <= sine_rom(3898);
     when "111100111011" => data <= sine_rom(3899);
     when "111100111100" => data <= sine_rom(3900);
     when "111100111101" => data <= sine_rom(3901);
     when "111100111110" => data <= sine_rom(3902);
     when "111100111111" => data <= sine_rom(3903);
     when "111101000000" => data <= sine_rom(3904);
     when "111101000001" => data <= sine_rom(3905);
     when "111101000010" => data <= sine_rom(3906);
     when "111101000011" => data <= sine_rom(3907);
     when "111101000100" => data <= sine_rom(3908);
     when "111101000101" => data <= sine_rom(3909);
     when "111101000110" => data <= sine_rom(3910);
     when "111101000111" => data <= sine_rom(3911);
     when "111101001000" => data <= sine_rom(3912);
     when "111101001001" => data <= sine_rom(3913);
     when "111101001010" => data <= sine_rom(3914);
     when "111101001011" => data <= sine_rom(3915);
     when "111101001100" => data <= sine_rom(3916);
     when "111101001101" => data <= sine_rom(3917);
     when "111101001110" => data <= sine_rom(3918);
     when "111101001111" => data <= sine_rom(3919);
     when "111101010000" => data <= sine_rom(3920);
     when "111101010001" => data <= sine_rom(3921);
     when "111101010010" => data <= sine_rom(3922);
     when "111101010011" => data <= sine_rom(3923);
     when "111101010100" => data <= sine_rom(3924);
     when "111101010101" => data <= sine_rom(3925);
     when "111101010110" => data <= sine_rom(3926);
     when "111101010111" => data <= sine_rom(3927);
     when "111101011000" => data <= sine_rom(3928);
     when "111101011001" => data <= sine_rom(3929);
     when "111101011010" => data <= sine_rom(3930);
     when "111101011011" => data <= sine_rom(3931);
     when "111101011100" => data <= sine_rom(3932);
     when "111101011101" => data <= sine_rom(3933);
     when "111101011110" => data <= sine_rom(3934);
     when "111101011111" => data <= sine_rom(3935);
     when "111101100000" => data <= sine_rom(3936);
     when "111101100001" => data <= sine_rom(3937);
     when "111101100010" => data <= sine_rom(3938);
     when "111101100011" => data <= sine_rom(3939);
     when "111101100100" => data <= sine_rom(3940);
     when "111101100101" => data <= sine_rom(3941);
     when "111101100110" => data <= sine_rom(3942);
     when "111101100111" => data <= sine_rom(3943);
     when "111101101000" => data <= sine_rom(3944);
     when "111101101001" => data <= sine_rom(3945);
     when "111101101010" => data <= sine_rom(3946);
     when "111101101011" => data <= sine_rom(3947);
     when "111101101100" => data <= sine_rom(3948);
     when "111101101101" => data <= sine_rom(3949);
     when "111101101110" => data <= sine_rom(3950);
     when "111101101111" => data <= sine_rom(3951);
     when "111101110000" => data <= sine_rom(3952);
     when "111101110001" => data <= sine_rom(3953);
     when "111101110010" => data <= sine_rom(3954);
     when "111101110011" => data <= sine_rom(3955);
     when "111101110100" => data <= sine_rom(3956);
     when "111101110101" => data <= sine_rom(3957);
     when "111101110110" => data <= sine_rom(3958);
     when "111101110111" => data <= sine_rom(3959);
     when "111101111000" => data <= sine_rom(3960);
     when "111101111001" => data <= sine_rom(3961);
     when "111101111010" => data <= sine_rom(3962);
     when "111101111011" => data <= sine_rom(3963);
     when "111101111100" => data <= sine_rom(3964);
     when "111101111101" => data <= sine_rom(3965);
     when "111101111110" => data <= sine_rom(3966);
     when "111101111111" => data <= sine_rom(3967);
     when "111110000000" => data <= sine_rom(3968);
     when "111110000001" => data <= sine_rom(3969);
     when "111110000010" => data <= sine_rom(3970);
     when "111110000011" => data <= sine_rom(3971);
     when "111110000100" => data <= sine_rom(3972);
     when "111110000101" => data <= sine_rom(3973);
     when "111110000110" => data <= sine_rom(3974);
     when "111110000111" => data <= sine_rom(3975);
     when "111110001000" => data <= sine_rom(3976);
     when "111110001001" => data <= sine_rom(3977);
     when "111110001010" => data <= sine_rom(3978);
     when "111110001011" => data <= sine_rom(3979);
     when "111110001100" => data <= sine_rom(3980);
     when "111110001101" => data <= sine_rom(3981);
     when "111110001110" => data <= sine_rom(3982);
     when "111110001111" => data <= sine_rom(3983);
     when "111110010000" => data <= sine_rom(3984);
     when "111110010001" => data <= sine_rom(3985);
     when "111110010010" => data <= sine_rom(3986);
     when "111110010011" => data <= sine_rom(3987);
     when "111110010100" => data <= sine_rom(3988);
     when "111110010101" => data <= sine_rom(3989);
     when "111110010110" => data <= sine_rom(3990);
     when "111110010111" => data <= sine_rom(3991);
     when "111110011000" => data <= sine_rom(3992);
     when "111110011001" => data <= sine_rom(3993);
     when "111110011010" => data <= sine_rom(3994);
     when "111110011011" => data <= sine_rom(3995);
     when "111110011100" => data <= sine_rom(3996);
     when "111110011101" => data <= sine_rom(3997);
     when "111110011110" => data <= sine_rom(3998);
     when "111110011111" => data <= sine_rom(3999);
     when "111110100000" => data <= sine_rom(4000);
     when "111110100001" => data <= sine_rom(4001);
     when "111110100010" => data <= sine_rom(4002);
     when "111110100011" => data <= sine_rom(4003);
     when "111110100100" => data <= sine_rom(4004);
     when "111110100101" => data <= sine_rom(4005);
     when "111110100110" => data <= sine_rom(4006);
     when "111110100111" => data <= sine_rom(4007);
     when "111110101000" => data <= sine_rom(4008);
     when "111110101001" => data <= sine_rom(4009);
     when "111110101010" => data <= sine_rom(4010);
     when "111110101011" => data <= sine_rom(4011);
     when "111110101100" => data <= sine_rom(4012);
     when "111110101101" => data <= sine_rom(4013);
     when "111110101110" => data <= sine_rom(4014);
     when "111110101111" => data <= sine_rom(4015);
     when "111110110000" => data <= sine_rom(4016);
     when "111110110001" => data <= sine_rom(4017);
     when "111110110010" => data <= sine_rom(4018);
     when "111110110011" => data <= sine_rom(4019);
     when "111110110100" => data <= sine_rom(4020);
     when "111110110101" => data <= sine_rom(4021);
     when "111110110110" => data <= sine_rom(4022);
     when "111110110111" => data <= sine_rom(4023);
     when "111110111000" => data <= sine_rom(4024);
     when "111110111001" => data <= sine_rom(4025);
     when "111110111010" => data <= sine_rom(4026);
     when "111110111011" => data <= sine_rom(4027);
     when "111110111100" => data <= sine_rom(4028);
     when "111110111101" => data <= sine_rom(4029);
     when "111110111110" => data <= sine_rom(4030);
     when "111110111111" => data <= sine_rom(4031);
     when "111111000000" => data <= sine_rom(4032);
     when "111111000001" => data <= sine_rom(4033);
     when "111111000010" => data <= sine_rom(4034);
     when "111111000011" => data <= sine_rom(4035);
     when "111111000100" => data <= sine_rom(4036);
     when "111111000101" => data <= sine_rom(4037);
     when "111111000110" => data <= sine_rom(4038);
     when "111111000111" => data <= sine_rom(4039);
     when "111111001000" => data <= sine_rom(4040);
     when "111111001001" => data <= sine_rom(4041);
     when "111111001010" => data <= sine_rom(4042);
     when "111111001011" => data <= sine_rom(4043);
     when "111111001100" => data <= sine_rom(4044);
     when "111111001101" => data <= sine_rom(4045);
     when "111111001110" => data <= sine_rom(4046);
     when "111111001111" => data <= sine_rom(4047);
     when "111111010000" => data <= sine_rom(4048);
     when "111111010001" => data <= sine_rom(4049);
     when "111111010010" => data <= sine_rom(4050);
     when "111111010011" => data <= sine_rom(4051);
     when "111111010100" => data <= sine_rom(4052);
     when "111111010101" => data <= sine_rom(4053);
     when "111111010110" => data <= sine_rom(4054);
     when "111111010111" => data <= sine_rom(4055);
     when "111111011000" => data <= sine_rom(4056);
     when "111111011001" => data <= sine_rom(4057);
     when "111111011010" => data <= sine_rom(4058);
     when "111111011011" => data <= sine_rom(4059);
     when "111111011100" => data <= sine_rom(4060);
     when "111111011101" => data <= sine_rom(4061);
     when "111111011110" => data <= sine_rom(4062);
     when "111111011111" => data <= sine_rom(4063);
     when "111111100000" => data <= sine_rom(4064);
     when "111111100001" => data <= sine_rom(4065);
     when "111111100010" => data <= sine_rom(4066);
     when "111111100011" => data <= sine_rom(4067);
     when "111111100100" => data <= sine_rom(4068);
     when "111111100101" => data <= sine_rom(4069);
     when "111111100110" => data <= sine_rom(4070);
     when "111111100111" => data <= sine_rom(4071);
     when "111111101000" => data <= sine_rom(4072);
     when "111111101001" => data <= sine_rom(4073);
     when "111111101010" => data <= sine_rom(4074);
     when "111111101011" => data <= sine_rom(4075);
     when "111111101100" => data <= sine_rom(4076);
     when "111111101101" => data <= sine_rom(4077);
     when "111111101110" => data <= sine_rom(4078);
     when "111111101111" => data <= sine_rom(4079);
     when "111111110000" => data <= sine_rom(4080);
     when "111111110001" => data <= sine_rom(4081);
     when "111111110010" => data <= sine_rom(4082);
     when "111111110011" => data <= sine_rom(4083);
     when "111111110100" => data <= sine_rom(4084);
     when "111111110101" => data <= sine_rom(4085);
     when "111111110110" => data <= sine_rom(4086);
     when "111111110111" => data <= sine_rom(4087);
     when "111111111000" => data <= sine_rom(4088);
     when "111111111001" => data <= sine_rom(4089);
     when "111111111010" => data <= sine_rom(4090);
     when "111111111011" => data <= sine_rom(4091);
     when "111111111100" => data <= sine_rom(4092);
     when "111111111101" => data <= sine_rom(4093);
     when "111111111110" => data <= sine_rom(4094);
     when "111111111111" => data <= sine_rom(4095);
     when others => data <= "000000000000";
    end case;
 end process;
end arch_Sine_LUT;
