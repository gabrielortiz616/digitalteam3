-------------------------------------------------------
--! @file
--! @brief Translate MIDI Note to phase increment sizer for the numerically controlled oscillator
-------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

--! Receive the MIDI Note number and returns the phase increment for the NCO
ENTITY MIDI_Increment_LUT IS
 port ( address : in std_logic_vector(7 downto 0); --! MIDI Note number
    data : out std_logic_vector(20 downto 0)); --! Phase increment size for NCO
 end entity MIDI_Increment_LUT;
 
--! Translate MIDI Note to phase increment sizer for the numerically controlled oscillator
 architecture arch_MIDI_Increment_LUT of MIDI_Increment_LUT is
    type mem is array ( 0 to 82) of std_logic_vector(20 downto 0);
    constant MIDI_rom : mem := (
    0 => "000000000010110100010", -- 1442 
    1 => "000000000010111111000", -- 1528 
    2 => "000000000011001010010", -- 1618 
    3 => "000000000011010110011", -- 1715 
    4 => "000000000011100011001", -- 1817 
    5 => "000000000011110000101", -- 1925 
    6 => "000000000011111110111", -- 2039 
    7 => "000000000100001110000", -- 2160 
    8 => "000000000100011110001", -- 2289 
    9 => "000000000100101111001", -- 2425 
    10 => "000000000101000001001", -- 2569 
    11 => "000000000101010100010", -- 2722 
    12 => "000000000101101000100", -- 2884 
    13 => "000000000101111101111", -- 3055 
    14 => "000000000110010100101", -- 3237 
    15 => "000000000110101100101", -- 3429 
    16 => "000000000111000110001", -- 3633 
    17 => "000000000111100001001", -- 3849 
    18 => "000000000111111101110", -- 4078 
    19 => "000000001000011100000", -- 4320 
    20 => "000000001000111100001", -- 4577 
    21 => "000000001001011110010", -- 4850 
    22 => "000000001010000010010", -- 5138 
    23 => "000000001010101000011", -- 5443 
    24 => "000000001011010000111", -- 5767 
    25 => "000000001011111011110", -- 6110 
    26 => "000000001100101001001", -- 6473 
    27 => "000000001101011001010", -- 6858 
    28 => "000000001110001100010", -- 7266 
    29 => "000000001111000010010", -- 7698 
    30 => "000000001111111011100", -- 8156 
    31 => "000000010000111000001", -- 8641 
    32 => "000000010001111000011", -- 9155 
    33 => "000000010010111100011", -- 9699 
    34 => "000000010100000100100", -- 10276 
    35 => "000000010101010000111", -- 10887 
    36 => "000000010110100001110", -- 11534 
    37 => "000000010111110111100", -- 12220 
    38 => "000000011001010010011", -- 12947 
    39 => "000000011010110010101", -- 13717 
    40 => "000000011100011000100", -- 14532 
    41 => "000000011110000100100", -- 15396 
    42 => "000000011111110111000", -- 16312 
    43 => "000000100001110000010", -- 17282 
    44 => "000000100011110000110", -- 18310 
    45 => "000000100101111000110", -- 19398 
    46 => "000000101000001001000", -- 20552 
    47 => "000000101010100001110", -- 21774 
    48 => "000000101101000011101", -- 23069 
    49 => "000000101111101111000", -- 24440 
    50 => "000000110010100100110", -- 25894 
    51 => "000000110101100101001", -- 27433 
    52 => "000000111000110001001", -- 29065 
    53 => "000000111100001001001", -- 30793 
    54 => "000000111111101110000", -- 32624 
    55 => "000001000011100000100", -- 34564 
    56 => "000001000111100001011", -- 36619 
    57 => "000001001011110001101", -- 38797 
    58 => "000001010000010010000", -- 41104 
    59 => "000001010101000011100", -- 43548 
    60 => "000001011010000111001", -- 46137 
    61 => "000001011111011110001", -- 48881 
    62 => "000001100101001001011", -- 51787 
    63 => "000001101011001010011", -- 54867 
    64 => "000001110001100010001", -- 58129 
    65 => "000001111000010010010", -- 61586 
    66 => "000001111111011100000", -- 65248 
    67 => "000010000111000001000", -- 69128 
    68 => "000010001111000010110", -- 73238 
    69 => "000010010111100011001", -- 77593 
    70 => "000010100000100011111", -- 82207 
    71 => "000010101010000111000", -- 87096 
    72 => "000010110100001110011", -- 92275 
    73 => "000010111110111100010", -- 97762 
    74 => "000011001010010010111", -- 103575 
    75 => "000011010110010100110", -- 109734 
    76 => "000011100011000100011", -- 116259 
    77 => "000011110000100100100", -- 123172 
    78 => "000011111110111000000", -- 130496 
    79 => "000100001110000010000", -- 138256 
    80 => "000100011110000101101", -- 146477 
    81 => "000100101111000110011", -- 155187 
    82 => "000101000001000111111"); -- 164415 
begin
 process (address)
 begin
  case address is
     when "00010101" => data <= MIDI_rom(0);  -- note 21
     when "00010110" => data <= MIDI_rom(1);  -- note 22
     when "00010111" => data <= MIDI_rom(2);  -- note 23
     when "00011000" => data <= MIDI_rom(3);  -- note 24
     when "00011001" => data <= MIDI_rom(4);  -- note 25
     when "00011010" => data <= MIDI_rom(5);  -- note 26
     when "00011011" => data <= MIDI_rom(6);  -- note 27
     when "00011100" => data <= MIDI_rom(7);  -- note 28
     when "00011101" => data <= MIDI_rom(8);  -- note 29
     when "00011110" => data <= MIDI_rom(9);  -- note 30
     when "00011111" => data <= MIDI_rom(10);  -- note 31
     when "00100000" => data <= MIDI_rom(11);  -- note 32
     when "00100001" => data <= MIDI_rom(12);  -- note 33
     when "00100010" => data <= MIDI_rom(13);  -- note 34
     when "00100011" => data <= MIDI_rom(14);  -- note 35
     when "00100100" => data <= MIDI_rom(15);  -- note 36
     when "00100101" => data <= MIDI_rom(16);  -- note 37
     when "00100110" => data <= MIDI_rom(17);  -- note 38
     when "00100111" => data <= MIDI_rom(18);  -- note 39
     when "00101000" => data <= MIDI_rom(19);  -- note 40
     when "00101001" => data <= MIDI_rom(20);  -- note 41
     when "00101010" => data <= MIDI_rom(21);  -- note 42
     when "00101011" => data <= MIDI_rom(22);  -- note 43
     when "00101100" => data <= MIDI_rom(23);  -- note 44
     when "00101101" => data <= MIDI_rom(24);  -- note 45
     when "00101110" => data <= MIDI_rom(25);  -- note 46
     when "00101111" => data <= MIDI_rom(26);  -- note 47
     when "00110000" => data <= MIDI_rom(27);  -- note 48
     when "00110001" => data <= MIDI_rom(28);  -- note 49
     when "00110010" => data <= MIDI_rom(29);  -- note 50
     when "00110011" => data <= MIDI_rom(30);  -- note 51
     when "00110100" => data <= MIDI_rom(31);  -- note 52
     when "00110101" => data <= MIDI_rom(32);  -- note 53
     when "00110110" => data <= MIDI_rom(33);  -- note 54
     when "00110111" => data <= MIDI_rom(34);  -- note 55
     when "00111000" => data <= MIDI_rom(35);  -- note 56
     when "00111001" => data <= MIDI_rom(36);  -- note 57
     when "00111010" => data <= MIDI_rom(37);  -- note 58
     when "00111011" => data <= MIDI_rom(38);  -- note 59
     when "00111100" => data <= MIDI_rom(39);  -- note 60
     when "00111101" => data <= MIDI_rom(40);  -- note 61
     when "00111110" => data <= MIDI_rom(41);  -- note 62
     when "00111111" => data <= MIDI_rom(42);  -- note 63
     when "01000000" => data <= MIDI_rom(43);  -- note 64
     when "01000001" => data <= MIDI_rom(44);  -- note 65
     when "01000010" => data <= MIDI_rom(45);  -- note 66
     when "01000011" => data <= MIDI_rom(46);  -- note 67
     when "01000100" => data <= MIDI_rom(47);  -- note 68
     when "01000101" => data <= MIDI_rom(48);  -- note 69
     when "01000110" => data <= MIDI_rom(49);  -- note 70
     when "01000111" => data <= MIDI_rom(50);  -- note 71
     when "01001000" => data <= MIDI_rom(51);  -- note 72
     when "01001001" => data <= MIDI_rom(52);  -- note 73
     when "01001010" => data <= MIDI_rom(53);  -- note 74
     when "01001011" => data <= MIDI_rom(54);  -- note 75
     when "01001100" => data <= MIDI_rom(55);  -- note 76
     when "01001101" => data <= MIDI_rom(56);  -- note 77
     when "01001110" => data <= MIDI_rom(57);  -- note 78
     when "01001111" => data <= MIDI_rom(58);  -- note 79
     when "01010000" => data <= MIDI_rom(59);  -- note 80
     when "01010001" => data <= MIDI_rom(60);  -- note 81
     when "01010010" => data <= MIDI_rom(61);  -- note 82
     when "01010011" => data <= MIDI_rom(62);  -- note 83
     when "01010100" => data <= MIDI_rom(63);  -- note 84
     when "01010101" => data <= MIDI_rom(64);  -- note 85
     when "01010110" => data <= MIDI_rom(65);  -- note 86
     when "01010111" => data <= MIDI_rom(66);  -- note 87
     when "01011000" => data <= MIDI_rom(67);  -- note 88
     when "01011001" => data <= MIDI_rom(68);  -- note 89
     when "01011010" => data <= MIDI_rom(69);  -- note 90
     when "01011011" => data <= MIDI_rom(70);  -- note 91
     when "01011100" => data <= MIDI_rom(71);  -- note 92
     when "01011101" => data <= MIDI_rom(72);  -- note 93
     when "01011110" => data <= MIDI_rom(73);  -- note 94
     when "01011111" => data <= MIDI_rom(74);  -- note 95
     when "01100000" => data <= MIDI_rom(75);  -- note 96
     when "01100001" => data <= MIDI_rom(76);  -- note 97
     when "01100010" => data <= MIDI_rom(77);  -- note 98
     when "01100011" => data <= MIDI_rom(78);  -- note 99
     when "01100100" => data <= MIDI_rom(79);  -- note 100
     when "01100101" => data <= MIDI_rom(80);  -- note 101
     when "01100110" => data <= MIDI_rom(81);  -- note 102
     when "01100111" => data <= MIDI_rom(82);  -- note 103
     when others => data <= "000000000000000000000";
    end case;
 end process;
end arch_MIDI_Increment_LUT;

