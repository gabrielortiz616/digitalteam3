LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.numeric_std.ALL;

ENTITY Square_DC_Reg IS
PORT(D : IN STD_LOGIC_VECTOR(6 DOWNTO 0); -- d_temputy cycle input.
     counter_size : IN STD_LOGIC_VECTOR(11 DOWNTO 0); -- counter size input.
	 reset : IN STD_LOGIC; -- Reset
	 clk : IN STD_LOGIC; -- clock.
	 slowclk : IN STD_LOGIC; -- clock.
	 Q : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)); -- output.
END Square_DC_Reg;

ARCHITECTURE arch_Square_DC_Reg OF Square_DC_Reg IS
signal d_temp: STD_LOGIC_VECTOR(6 DOWNTO 0) :="1000010"; -- d_temputy cycle input.
BEGIN
    PROCESS(clk, reset)
    BEGIN
	d_temp <= D;
        IF reset = '0' THEN
				Q <= (others => '0');
        ELSIF rising_edge(clk) THEN
            IF slowclk ='1' THEN
                IF d_temp >= "0000000" AND d_temp<"0000010" THEN
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7))); 
			    ELSIF d_temp >= "0000010" AND d_temp<"0000011" THEN
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));      
                ELSIF d_temp >= "0000011" AND d_temp<"0000100" THEN
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));                     
                ELSIF d_temp >= "0000100" AND d_temp<"0000101" THEN
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));					 
                ELSIF d_temp >= "0000101" AND d_temp<"0000110" THEN
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0000110" AND d_temp<"0000111" THEN
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6)));                
			    ELSIF d_temp >= "0000111" AND d_temp<"0001000" THEN
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0001000" AND d_temp<"0001001" THEN                        
 					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4)));
                ELSIF d_temp >= "0001001" AND d_temp<"0001010" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0001010" AND d_temp<"0001011" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));
                ELSIF d_temp >= "0001011" AND d_temp<"0001100" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                ELSIF d_temp >= "0001100" AND d_temp<"0001101" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5)));                                     
                ELSIF d_temp >= "0001101" AND d_temp<"0001110" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                ELSIF d_temp >= "0001110" AND d_temp<"0001111" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6)));
                ELSIF d_temp >= "0001111" AND d_temp<"0010000" THEN                        
 					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0010000" AND d_temp<"0010001" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3)));
                ELSIF d_temp >= "0010001" AND d_temp<"0010010" THEN                        
 					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7))); 
                ELSIF d_temp >= "0010010" AND d_temp<"0010011" THEN                        
 					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6)));  
                ELSIF d_temp >= "0010011" AND d_temp<"0010100" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0010100" AND d_temp<"0010101" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));
                ELSIF d_temp >= "0010101" AND d_temp<"0010110" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0010110" AND d_temp<"0010111" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))); 
                ELSIF d_temp >= "0010111" AND d_temp<"0011000" THEN                        
    				 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0011000" AND d_temp<"0011001" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4)));      
                ELSIF d_temp >= "0011001" AND d_temp<"0011010" THEN                        
					 Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                ELSIF d_temp >= "0011010" AND d_temp<"0011011" THEN                        
                     Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));  
                ELSIF d_temp >= "0011011" AND d_temp<"0011100" THEN                        
                     Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                ELSIF d_temp >= "0011100" AND d_temp<"0011101" THEN                        
                     Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5)));  
                ELSIF d_temp >= "0011101" AND d_temp<"0011110" THEN                        
                     Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                ELSIF d_temp >= "0011110" AND d_temp<"0011111" THEN                         
                     Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 6)));   
                ELSIF d_temp >= "0100000" AND d_temp<"0100001" THEN                         
                     Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 7)));                                            
                ELSIF d_temp >= "0100001" AND d_temp<"0100010" THEN                         
                     Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)));  
                ELSIF d_temp >= "0100010" AND d_temp<"0100011" THEN
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7))); 
                 ELSIF d_temp >= "0100011" AND d_temp<"0100100" THEN
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));      
                 ELSIF d_temp >= "0100100" AND d_temp<"0100101" THEN
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));                     
                 ELSIF d_temp >= "0100101" AND d_temp<"0100110" THEN
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));                     
                 ELSIF d_temp >= "0100110" AND d_temp<"0100111" THEN
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "0100111" AND d_temp<"0101000" THEN
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6)));                
                 ELSIF d_temp >= "0101000" AND d_temp<"0101001" THEN
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "0101001" AND d_temp<"0101010" THEN                        
                       Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4)));
                 ELSIF d_temp >= "0101010" AND d_temp<"0101011" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "0101011" AND d_temp<"0101100" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));
                 ELSIF d_temp >= "0101100" AND d_temp<"0101101" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                 ELSIF d_temp >= "0101101" AND d_temp<"0101110" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5)));                                     
                 ELSIF d_temp >= "0101110" AND d_temp<"0101111" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                 ELSIF d_temp >= "0101111" AND d_temp<"0110000" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6)));
                 ELSIF d_temp >= "0110000" AND d_temp<"0110001" THEN                        
                       Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "0110001" AND d_temp<"0110010" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 3)));
                 ELSIF d_temp >= "0110010" AND d_temp<"0110011" THEN                        
                       Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7))); 
                 ELSIF d_temp >= "0110011" AND d_temp<"0110100" THEN                        
                       Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6)));  
                 ELSIF d_temp >= "0110100" AND d_temp<"0110101" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "0110101" AND d_temp<"0110110" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));
                 ELSIF d_temp >= "0110110" AND d_temp<"0110111" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "0110111" AND d_temp<"0111000" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))); 
                 ELSIF d_temp >= "0111000" AND d_temp<"0111001" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "0111001" AND d_temp<"0111010" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 4)));      
                 ELSIF d_temp >= "0111010" AND d_temp<"0111011" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                 ELSIF d_temp >= "0111100" AND d_temp<"0111101" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));  
                 ELSIF d_temp >= "0111101" AND d_temp<"0111110" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                 ELSIF d_temp >= "0111110" AND d_temp<"0111111" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 5)));  
                 ELSIF d_temp >= "0111111" AND d_temp<"1000000" THEN                        
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                 ELSIF d_temp >= "1000000" AND d_temp<"1000001" THEN                         
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)) + unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 6)));   
                 ELSIF d_temp >= "1000001" AND d_temp<"1000010" THEN                         
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1))+ unsigned(shift_right(unsigned(counter_size), 7)));                                            
                 ELSIF d_temp >= "1000010" AND d_temp<"1000011" THEN                         
                      Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 1)));     
                      ELSIF d_temp >= "1000011" AND d_temp<"1000100" THEN
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));                     
                      ELSIF d_temp >= "1000100" AND d_temp<"1000101" THEN
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));                     
                      ELSIF d_temp >= "1000101" AND d_temp<"1000110" THEN
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1000110" AND d_temp<"1000111" THEN
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6)));                
                      ELSIF d_temp >= "1000111" AND d_temp<"1001000" THEN
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1001000" AND d_temp<"1001001" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4)));
                      ELSIF d_temp >= "1001001" AND d_temp<"1001010" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1001010" AND d_temp<"1001011" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));
                      ELSIF d_temp >= "1001011" AND d_temp<"1001100" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                      ELSIF d_temp >= "1001100" AND d_temp<"1001101" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5)));                                     
                      ELSIF d_temp >= "1001101" AND d_temp<"1001110" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                      ELSIF d_temp >= "1001110" AND d_temp<"1001111" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6)));
                      ELSIF d_temp >= "1001111" AND d_temp<"1010000" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1010000" AND d_temp<"1010001" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 3)));
                      ELSIF d_temp >= "1010001" AND d_temp<"1010010" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7))); 
                      ELSIF d_temp >= "1010010" AND d_temp<"1010011" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6)));  
                      ELSIF d_temp >= "1010011" AND d_temp<"1010100" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1010100" AND d_temp<"1010101" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));
                      ELSIF d_temp >= "1010101" AND d_temp<"1010110" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1010110" AND d_temp<"1010111" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))); 
                      ELSIF d_temp >= "1010111" AND d_temp<"1011000" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1011000" AND d_temp<"1011001" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 4)));      
                      ELSIF d_temp >= "1011001" AND d_temp<"1011010" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                      ELSIF d_temp >= "1011010" AND d_temp<"1011011" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));  
                      ELSIF d_temp >= "1011011" AND d_temp<"1011100" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                      ELSIF d_temp >= "1011100" AND d_temp<"1011101" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 5)));  
                      ELSIF d_temp >= "1011101" AND d_temp<"1011110" THEN                        
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                      ELSIF d_temp >= "1011110" AND d_temp<"1011111" THEN                         
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 6)));   
                      ELSIF d_temp >= "1100000" AND d_temp<"1100001" THEN                         
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)) + unsigned(shift_right(unsigned(counter_size), 7)));                                            
                      ELSIF d_temp >= "1100001" AND d_temp<"1100010" THEN                         
                           Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 2)));  
                      ELSIF d_temp >= "1100010" AND d_temp<"1100011" THEN
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7))); 
                       ELSIF d_temp >= "1100011" AND d_temp<"1100100" THEN
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));      
                       ELSIF d_temp >= "1100100" AND d_temp<"1100101" THEN
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));                     
                       ELSIF d_temp >= "1100101" AND d_temp<"1100110" THEN
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));                     
                       ELSIF d_temp >= "1100110" AND d_temp<"1100111" THEN
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                       ELSIF d_temp >= "1100111" AND d_temp<"1101000" THEN
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6)));                
                       ELSIF d_temp >= "1101000" AND d_temp<"1101001" THEN
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                       ELSIF d_temp >= "1101001" AND d_temp<"1101010" THEN                        
                             Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 4)));
                       ELSIF d_temp >= "1101010" AND d_temp<"1101011" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                       ELSIF d_temp >= "1101011" AND d_temp<"1101100" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));
                       ELSIF d_temp >= "1101100" AND d_temp<"1101101" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                       ELSIF d_temp >= "1101101" AND d_temp<"1101110" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 5)));                                     
                       ELSIF d_temp >= "1101110" AND d_temp<"1101111" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                       ELSIF d_temp >= "1101111" AND d_temp<"1110000" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 6)));
                       ELSIF d_temp >= "1110000" AND d_temp<"1110001" THEN                        
                             Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3))+ unsigned(shift_right(unsigned(counter_size), 7)));
                       ELSIF d_temp >= "1110001" AND d_temp<"1110010" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 3)));
                       ELSIF d_temp >= "1110010" AND d_temp<"1110011" THEN                        
                             Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7))); 
                       ELSIF d_temp >= "1110011" AND d_temp<"1110100" THEN                        
                             Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 6)));  
                       ELSIF d_temp >= "1110100" AND d_temp<"1110101" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)) + unsigned(shift_right(unsigned(counter_size), 7)));
                       ELSIF d_temp >= "1110101" AND d_temp<"1110110" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 5)));
                       ELSIF d_temp >= "1110110" AND d_temp<"1110111" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));
                       ELSIF d_temp >= "1110111" AND d_temp<"1111000" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 6))); 
                       ELSIF d_temp >= "1111000" AND d_temp<"1111001" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4))+ unsigned(shift_right(unsigned(counter_size), 7)));
                       ELSIF d_temp >= "1111001" AND d_temp<"1111010" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 4)));      
                       ELSIF d_temp >= "1111010" AND d_temp<"1111011" THEN                        
                            Q <= std_logic_vector(  unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                       ELSIF d_temp >= "1111100" AND d_temp<"1111101" THEN                        
                            Q <= std_logic_vector( unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 6)));  
                       ELSIF d_temp >= "1111101" AND d_temp<"1111110" THEN                        
                            Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 5))+ unsigned(shift_right(unsigned(counter_size), 7)));  
                       ELSIF d_temp >= "1111110" AND d_temp<"1111111" THEN                        
                            Q <= std_logic_vector(unsigned(shift_right(unsigned(counter_size), 6)));  
                ELSE                     
                     Q <= std_logic_vector(shift_right(unsigned(counter_size), 1)); 
                END IF;                                                                                                        			         
			END IF;
        END IF;
    END PROCESS;
END arch_Square_DC_Reg;
