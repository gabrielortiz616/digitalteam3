library ieee;
use ieee.std_logic_1164.all;
entity Sawtooth_LUT is
 port ( address : in std_logic_vector(11 downto 0);
    data : out std_logic_vector(11 downto 0));
 end entity Sawtooth_LUT;
 architecture arch_Sawtooth_LUT of Sawtooth_LUT is
    type mem is array ( 0 to 2**12 - 1) of std_logic_vector(11 downto 0);
    constant saw_rom : mem := (
    0 => "000000000000",
    1 => "000000000001",
    2 => "000000000010",
    3 => "000000000011",
    4 => "000000000100",
    5 => "000000000101",
    6 => "000000000110",
    7 => "000000000111",
    8 => "000000001000",
    9 => "000000001001",
    10 => "000000001010",
    11 => "000000001011",
    12 => "000000001100",
    13 => "000000001101",
    14 => "000000001110",
    15 => "000000001111",
    16 => "000000010000",
    17 => "000000010001",
    18 => "000000010010",
    19 => "000000010011",
    20 => "000000010100",
    21 => "000000010101",
    22 => "000000010110",
    23 => "000000010111",
    24 => "000000011000",
    25 => "000000011001",
    26 => "000000011010",
    27 => "000000011011",
    28 => "000000011100",
    29 => "000000011101",
    30 => "000000011110",
    31 => "000000011111",
    32 => "000000100000",
    33 => "000000100001",
    34 => "000000100010",
    35 => "000000100011",
    36 => "000000100100",
    37 => "000000100101",
    38 => "000000100110",
    39 => "000000100111",
    40 => "000000101000",
    41 => "000000101001",
    42 => "000000101010",
    43 => "000000101011",
    44 => "000000101100",
    45 => "000000101101",
    46 => "000000101110",
    47 => "000000101111",
    48 => "000000110000",
    49 => "000000110001",
    50 => "000000110010",
    51 => "000000110011",
    52 => "000000110100",
    53 => "000000110101",
    54 => "000000110110",
    55 => "000000110111",
    56 => "000000111000",
    57 => "000000111001",
    58 => "000000111010",
    59 => "000000111011",
    60 => "000000111100",
    61 => "000000111101",
    62 => "000000111110",
    63 => "000000111111",
    64 => "000001000000",
    65 => "000001000001",
    66 => "000001000010",
    67 => "000001000011",
    68 => "000001000100",
    69 => "000001000101",
    70 => "000001000110",
    71 => "000001000111",
    72 => "000001001000",
    73 => "000001001001",
    74 => "000001001010",
    75 => "000001001011",
    76 => "000001001100",
    77 => "000001001101",
    78 => "000001001110",
    79 => "000001001111",
    80 => "000001010000",
    81 => "000001010001",
    82 => "000001010010",
    83 => "000001010011",
    84 => "000001010100",
    85 => "000001010101",
    86 => "000001010110",
    87 => "000001010111",
    88 => "000001011000",
    89 => "000001011001",
    90 => "000001011010",
    91 => "000001011011",
    92 => "000001011100",
    93 => "000001011101",
    94 => "000001011110",
    95 => "000001011111",
    96 => "000001100000",
    97 => "000001100001",
    98 => "000001100010",
    99 => "000001100011",
    100 => "000001100100",
    101 => "000001100101",
    102 => "000001100110",
    103 => "000001100111",
    104 => "000001101000",
    105 => "000001101001",
    106 => "000001101010",
    107 => "000001101011",
    108 => "000001101100",
    109 => "000001101101",
    110 => "000001101110",
    111 => "000001101111",
    112 => "000001110000",
    113 => "000001110001",
    114 => "000001110010",
    115 => "000001110011",
    116 => "000001110100",
    117 => "000001110101",
    118 => "000001110110",
    119 => "000001110111",
    120 => "000001111000",
    121 => "000001111001",
    122 => "000001111010",
    123 => "000001111011",
    124 => "000001111100",
    125 => "000001111101",
    126 => "000001111110",
    127 => "000001111111",
    128 => "000010000000",
    129 => "000010000001",
    130 => "000010000010",
    131 => "000010000011",
    132 => "000010000100",
    133 => "000010000101",
    134 => "000010000110",
    135 => "000010000111",
    136 => "000010001000",
    137 => "000010001001",
    138 => "000010001010",
    139 => "000010001011",
    140 => "000010001100",
    141 => "000010001101",
    142 => "000010001110",
    143 => "000010001111",
    144 => "000010010000",
    145 => "000010010001",
    146 => "000010010010",
    147 => "000010010011",
    148 => "000010010100",
    149 => "000010010101",
    150 => "000010010110",
    151 => "000010010111",
    152 => "000010011000",
    153 => "000010011001",
    154 => "000010011010",
    155 => "000010011011",
    156 => "000010011100",
    157 => "000010011101",
    158 => "000010011110",
    159 => "000010011111",
    160 => "000010100000",
    161 => "000010100001",
    162 => "000010100010",
    163 => "000010100011",
    164 => "000010100100",
    165 => "000010100101",
    166 => "000010100110",
    167 => "000010100111",
    168 => "000010101000",
    169 => "000010101001",
    170 => "000010101010",
    171 => "000010101011",
    172 => "000010101100",
    173 => "000010101101",
    174 => "000010101110",
    175 => "000010101111",
    176 => "000010110000",
    177 => "000010110001",
    178 => "000010110010",
    179 => "000010110011",
    180 => "000010110100",
    181 => "000010110101",
    182 => "000010110110",
    183 => "000010110111",
    184 => "000010111000",
    185 => "000010111001",
    186 => "000010111010",
    187 => "000010111011",
    188 => "000010111100",
    189 => "000010111101",
    190 => "000010111110",
    191 => "000010111111",
    192 => "000011000000",
    193 => "000011000001",
    194 => "000011000010",
    195 => "000011000011",
    196 => "000011000100",
    197 => "000011000101",
    198 => "000011000110",
    199 => "000011000111",
    200 => "000011001000",
    201 => "000011001001",
    202 => "000011001010",
    203 => "000011001011",
    204 => "000011001100",
    205 => "000011001101",
    206 => "000011001110",
    207 => "000011001111",
    208 => "000011010000",
    209 => "000011010001",
    210 => "000011010010",
    211 => "000011010011",
    212 => "000011010100",
    213 => "000011010101",
    214 => "000011010110",
    215 => "000011010111",
    216 => "000011011000",
    217 => "000011011001",
    218 => "000011011010",
    219 => "000011011011",
    220 => "000011011100",
    221 => "000011011101",
    222 => "000011011110",
    223 => "000011011111",
    224 => "000011100000",
    225 => "000011100001",
    226 => "000011100010",
    227 => "000011100011",
    228 => "000011100100",
    229 => "000011100101",
    230 => "000011100110",
    231 => "000011100111",
    232 => "000011101000",
    233 => "000011101001",
    234 => "000011101010",
    235 => "000011101011",
    236 => "000011101100",
    237 => "000011101101",
    238 => "000011101110",
    239 => "000011101111",
    240 => "000011110000",
    241 => "000011110001",
    242 => "000011110010",
    243 => "000011110011",
    244 => "000011110100",
    245 => "000011110101",
    246 => "000011110110",
    247 => "000011110111",
    248 => "000011111000",
    249 => "000011111001",
    250 => "000011111010",
    251 => "000011111011",
    252 => "000011111100",
    253 => "000011111101",
    254 => "000011111110",
    255 => "000011111111",
    256 => "000100000000",
    257 => "000100000001",
    258 => "000100000010",
    259 => "000100000011",
    260 => "000100000100",
    261 => "000100000101",
    262 => "000100000110",
    263 => "000100000111",
    264 => "000100001000",
    265 => "000100001001",
    266 => "000100001010",
    267 => "000100001011",
    268 => "000100001100",
    269 => "000100001101",
    270 => "000100001110",
    271 => "000100001111",
    272 => "000100010000",
    273 => "000100010001",
    274 => "000100010010",
    275 => "000100010011",
    276 => "000100010100",
    277 => "000100010101",
    278 => "000100010110",
    279 => "000100010111",
    280 => "000100011000",
    281 => "000100011001",
    282 => "000100011010",
    283 => "000100011011",
    284 => "000100011100",
    285 => "000100011101",
    286 => "000100011110",
    287 => "000100011111",
    288 => "000100100000",
    289 => "000100100001",
    290 => "000100100010",
    291 => "000100100011",
    292 => "000100100100",
    293 => "000100100101",
    294 => "000100100110",
    295 => "000100100111",
    296 => "000100101000",
    297 => "000100101001",
    298 => "000100101010",
    299 => "000100101011",
    300 => "000100101100",
    301 => "000100101101",
    302 => "000100101110",
    303 => "000100101111",
    304 => "000100110000",
    305 => "000100110001",
    306 => "000100110010",
    307 => "000100110011",
    308 => "000100110100",
    309 => "000100110101",
    310 => "000100110110",
    311 => "000100110111",
    312 => "000100111000",
    313 => "000100111001",
    314 => "000100111010",
    315 => "000100111011",
    316 => "000100111100",
    317 => "000100111101",
    318 => "000100111110",
    319 => "000100111111",
    320 => "000101000000",
    321 => "000101000001",
    322 => "000101000010",
    323 => "000101000011",
    324 => "000101000100",
    325 => "000101000101",
    326 => "000101000110",
    327 => "000101000111",
    328 => "000101001000",
    329 => "000101001001",
    330 => "000101001010",
    331 => "000101001011",
    332 => "000101001100",
    333 => "000101001101",
    334 => "000101001110",
    335 => "000101001111",
    336 => "000101010000",
    337 => "000101010001",
    338 => "000101010010",
    339 => "000101010011",
    340 => "000101010100",
    341 => "000101010101",
    342 => "000101010110",
    343 => "000101010111",
    344 => "000101011000",
    345 => "000101011001",
    346 => "000101011010",
    347 => "000101011011",
    348 => "000101011100",
    349 => "000101011101",
    350 => "000101011110",
    351 => "000101011111",
    352 => "000101100000",
    353 => "000101100001",
    354 => "000101100010",
    355 => "000101100011",
    356 => "000101100100",
    357 => "000101100101",
    358 => "000101100110",
    359 => "000101100111",
    360 => "000101101000",
    361 => "000101101001",
    362 => "000101101010",
    363 => "000101101011",
    364 => "000101101100",
    365 => "000101101101",
    366 => "000101101110",
    367 => "000101101111",
    368 => "000101110000",
    369 => "000101110001",
    370 => "000101110010",
    371 => "000101110011",
    372 => "000101110100",
    373 => "000101110101",
    374 => "000101110110",
    375 => "000101110111",
    376 => "000101111000",
    377 => "000101111001",
    378 => "000101111010",
    379 => "000101111011",
    380 => "000101111100",
    381 => "000101111101",
    382 => "000101111110",
    383 => "000101111111",
    384 => "000110000000",
    385 => "000110000001",
    386 => "000110000010",
    387 => "000110000011",
    388 => "000110000100",
    389 => "000110000101",
    390 => "000110000110",
    391 => "000110000111",
    392 => "000110001000",
    393 => "000110001001",
    394 => "000110001010",
    395 => "000110001011",
    396 => "000110001100",
    397 => "000110001101",
    398 => "000110001110",
    399 => "000110001111",
    400 => "000110010000",
    401 => "000110010001",
    402 => "000110010010",
    403 => "000110010011",
    404 => "000110010100",
    405 => "000110010101",
    406 => "000110010110",
    407 => "000110010111",
    408 => "000110011000",
    409 => "000110011001",
    410 => "000110011010",
    411 => "000110011011",
    412 => "000110011100",
    413 => "000110011101",
    414 => "000110011110",
    415 => "000110011111",
    416 => "000110100000",
    417 => "000110100001",
    418 => "000110100010",
    419 => "000110100011",
    420 => "000110100100",
    421 => "000110100101",
    422 => "000110100110",
    423 => "000110100111",
    424 => "000110101000",
    425 => "000110101001",
    426 => "000110101010",
    427 => "000110101011",
    428 => "000110101100",
    429 => "000110101101",
    430 => "000110101110",
    431 => "000110101111",
    432 => "000110110000",
    433 => "000110110001",
    434 => "000110110010",
    435 => "000110110011",
    436 => "000110110100",
    437 => "000110110101",
    438 => "000110110110",
    439 => "000110110111",
    440 => "000110111000",
    441 => "000110111001",
    442 => "000110111010",
    443 => "000110111011",
    444 => "000110111100",
    445 => "000110111101",
    446 => "000110111110",
    447 => "000110111111",
    448 => "000111000000",
    449 => "000111000001",
    450 => "000111000010",
    451 => "000111000011",
    452 => "000111000100",
    453 => "000111000101",
    454 => "000111000110",
    455 => "000111000111",
    456 => "000111001000",
    457 => "000111001001",
    458 => "000111001010",
    459 => "000111001011",
    460 => "000111001100",
    461 => "000111001101",
    462 => "000111001110",
    463 => "000111001111",
    464 => "000111010000",
    465 => "000111010001",
    466 => "000111010010",
    467 => "000111010011",
    468 => "000111010100",
    469 => "000111010101",
    470 => "000111010110",
    471 => "000111010111",
    472 => "000111011000",
    473 => "000111011001",
    474 => "000111011010",
    475 => "000111011011",
    476 => "000111011100",
    477 => "000111011101",
    478 => "000111011110",
    479 => "000111011111",
    480 => "000111100000",
    481 => "000111100001",
    482 => "000111100010",
    483 => "000111100011",
    484 => "000111100100",
    485 => "000111100101",
    486 => "000111100110",
    487 => "000111100111",
    488 => "000111101000",
    489 => "000111101001",
    490 => "000111101010",
    491 => "000111101011",
    492 => "000111101100",
    493 => "000111101101",
    494 => "000111101110",
    495 => "000111101111",
    496 => "000111110000",
    497 => "000111110001",
    498 => "000111110010",
    499 => "000111110011",
    500 => "000111110100",
    501 => "000111110101",
    502 => "000111110110",
    503 => "000111110111",
    504 => "000111111000",
    505 => "000111111001",
    506 => "000111111010",
    507 => "000111111011",
    508 => "000111111100",
    509 => "000111111101",
    510 => "000111111110",
    511 => "000111111111",
    512 => "001000000000",
    513 => "001000000001",
    514 => "001000000010",
    515 => "001000000011",
    516 => "001000000100",
    517 => "001000000101",
    518 => "001000000110",
    519 => "001000000111",
    520 => "001000001000",
    521 => "001000001001",
    522 => "001000001010",
    523 => "001000001011",
    524 => "001000001100",
    525 => "001000001101",
    526 => "001000001110",
    527 => "001000001111",
    528 => "001000010000",
    529 => "001000010001",
    530 => "001000010010",
    531 => "001000010011",
    532 => "001000010100",
    533 => "001000010101",
    534 => "001000010110",
    535 => "001000010111",
    536 => "001000011000",
    537 => "001000011001",
    538 => "001000011010",
    539 => "001000011011",
    540 => "001000011100",
    541 => "001000011101",
    542 => "001000011110",
    543 => "001000011111",
    544 => "001000100000",
    545 => "001000100001",
    546 => "001000100010",
    547 => "001000100011",
    548 => "001000100100",
    549 => "001000100101",
    550 => "001000100110",
    551 => "001000100111",
    552 => "001000101000",
    553 => "001000101001",
    554 => "001000101010",
    555 => "001000101011",
    556 => "001000101100",
    557 => "001000101101",
    558 => "001000101110",
    559 => "001000101111",
    560 => "001000110000",
    561 => "001000110001",
    562 => "001000110010",
    563 => "001000110011",
    564 => "001000110100",
    565 => "001000110101",
    566 => "001000110110",
    567 => "001000110111",
    568 => "001000111000",
    569 => "001000111001",
    570 => "001000111010",
    571 => "001000111011",
    572 => "001000111100",
    573 => "001000111101",
    574 => "001000111110",
    575 => "001000111111",
    576 => "001001000000",
    577 => "001001000001",
    578 => "001001000010",
    579 => "001001000011",
    580 => "001001000100",
    581 => "001001000101",
    582 => "001001000110",
    583 => "001001000111",
    584 => "001001001000",
    585 => "001001001001",
    586 => "001001001010",
    587 => "001001001011",
    588 => "001001001100",
    589 => "001001001101",
    590 => "001001001110",
    591 => "001001001111",
    592 => "001001010000",
    593 => "001001010001",
    594 => "001001010010",
    595 => "001001010011",
    596 => "001001010100",
    597 => "001001010101",
    598 => "001001010110",
    599 => "001001010111",
    600 => "001001011000",
    601 => "001001011001",
    602 => "001001011010",
    603 => "001001011011",
    604 => "001001011100",
    605 => "001001011101",
    606 => "001001011110",
    607 => "001001011111",
    608 => "001001100000",
    609 => "001001100001",
    610 => "001001100010",
    611 => "001001100011",
    612 => "001001100100",
    613 => "001001100101",
    614 => "001001100110",
    615 => "001001100111",
    616 => "001001101000",
    617 => "001001101001",
    618 => "001001101010",
    619 => "001001101011",
    620 => "001001101100",
    621 => "001001101101",
    622 => "001001101110",
    623 => "001001101111",
    624 => "001001110000",
    625 => "001001110001",
    626 => "001001110010",
    627 => "001001110011",
    628 => "001001110100",
    629 => "001001110101",
    630 => "001001110110",
    631 => "001001110111",
    632 => "001001111000",
    633 => "001001111001",
    634 => "001001111010",
    635 => "001001111011",
    636 => "001001111100",
    637 => "001001111101",
    638 => "001001111110",
    639 => "001001111111",
    640 => "001010000000",
    641 => "001010000001",
    642 => "001010000010",
    643 => "001010000011",
    644 => "001010000100",
    645 => "001010000101",
    646 => "001010000110",
    647 => "001010000111",
    648 => "001010001000",
    649 => "001010001001",
    650 => "001010001010",
    651 => "001010001011",
    652 => "001010001100",
    653 => "001010001101",
    654 => "001010001110",
    655 => "001010001111",
    656 => "001010010000",
    657 => "001010010001",
    658 => "001010010010",
    659 => "001010010011",
    660 => "001010010100",
    661 => "001010010101",
    662 => "001010010110",
    663 => "001010010111",
    664 => "001010011000",
    665 => "001010011001",
    666 => "001010011010",
    667 => "001010011011",
    668 => "001010011100",
    669 => "001010011101",
    670 => "001010011110",
    671 => "001010011111",
    672 => "001010100000",
    673 => "001010100001",
    674 => "001010100010",
    675 => "001010100011",
    676 => "001010100100",
    677 => "001010100101",
    678 => "001010100110",
    679 => "001010100111",
    680 => "001010101000",
    681 => "001010101001",
    682 => "001010101010",
    683 => "001010101011",
    684 => "001010101100",
    685 => "001010101101",
    686 => "001010101110",
    687 => "001010101111",
    688 => "001010110000",
    689 => "001010110001",
    690 => "001010110010",
    691 => "001010110011",
    692 => "001010110100",
    693 => "001010110101",
    694 => "001010110110",
    695 => "001010110111",
    696 => "001010111000",
    697 => "001010111001",
    698 => "001010111010",
    699 => "001010111011",
    700 => "001010111100",
    701 => "001010111101",
    702 => "001010111110",
    703 => "001010111111",
    704 => "001011000000",
    705 => "001011000001",
    706 => "001011000010",
    707 => "001011000011",
    708 => "001011000100",
    709 => "001011000101",
    710 => "001011000110",
    711 => "001011000111",
    712 => "001011001000",
    713 => "001011001001",
    714 => "001011001010",
    715 => "001011001011",
    716 => "001011001100",
    717 => "001011001101",
    718 => "001011001110",
    719 => "001011001111",
    720 => "001011010000",
    721 => "001011010001",
    722 => "001011010010",
    723 => "001011010011",
    724 => "001011010100",
    725 => "001011010101",
    726 => "001011010110",
    727 => "001011010111",
    728 => "001011011000",
    729 => "001011011001",
    730 => "001011011010",
    731 => "001011011011",
    732 => "001011011100",
    733 => "001011011101",
    734 => "001011011110",
    735 => "001011011111",
    736 => "001011100000",
    737 => "001011100001",
    738 => "001011100010",
    739 => "001011100011",
    740 => "001011100100",
    741 => "001011100101",
    742 => "001011100110",
    743 => "001011100111",
    744 => "001011101000",
    745 => "001011101001",
    746 => "001011101010",
    747 => "001011101011",
    748 => "001011101100",
    749 => "001011101101",
    750 => "001011101110",
    751 => "001011101111",
    752 => "001011110000",
    753 => "001011110001",
    754 => "001011110010",
    755 => "001011110011",
    756 => "001011110100",
    757 => "001011110101",
    758 => "001011110110",
    759 => "001011110111",
    760 => "001011111000",
    761 => "001011111001",
    762 => "001011111010",
    763 => "001011111011",
    764 => "001011111100",
    765 => "001011111101",
    766 => "001011111110",
    767 => "001011111111",
    768 => "001100000000",
    769 => "001100000001",
    770 => "001100000010",
    771 => "001100000011",
    772 => "001100000100",
    773 => "001100000101",
    774 => "001100000110",
    775 => "001100000111",
    776 => "001100001000",
    777 => "001100001001",
    778 => "001100001010",
    779 => "001100001011",
    780 => "001100001100",
    781 => "001100001101",
    782 => "001100001110",
    783 => "001100001111",
    784 => "001100010000",
    785 => "001100010001",
    786 => "001100010010",
    787 => "001100010011",
    788 => "001100010100",
    789 => "001100010101",
    790 => "001100010110",
    791 => "001100010111",
    792 => "001100011000",
    793 => "001100011001",
    794 => "001100011010",
    795 => "001100011011",
    796 => "001100011100",
    797 => "001100011101",
    798 => "001100011110",
    799 => "001100011111",
    800 => "001100100000",
    801 => "001100100001",
    802 => "001100100010",
    803 => "001100100011",
    804 => "001100100100",
    805 => "001100100101",
    806 => "001100100110",
    807 => "001100100111",
    808 => "001100101000",
    809 => "001100101001",
    810 => "001100101010",
    811 => "001100101011",
    812 => "001100101100",
    813 => "001100101101",
    814 => "001100101110",
    815 => "001100101111",
    816 => "001100110000",
    817 => "001100110001",
    818 => "001100110010",
    819 => "001100110011",
    820 => "001100110100",
    821 => "001100110101",
    822 => "001100110110",
    823 => "001100110111",
    824 => "001100111000",
    825 => "001100111001",
    826 => "001100111010",
    827 => "001100111011",
    828 => "001100111100",
    829 => "001100111101",
    830 => "001100111110",
    831 => "001100111111",
    832 => "001101000000",
    833 => "001101000001",
    834 => "001101000010",
    835 => "001101000011",
    836 => "001101000100",
    837 => "001101000101",
    838 => "001101000110",
    839 => "001101000111",
    840 => "001101001000",
    841 => "001101001001",
    842 => "001101001010",
    843 => "001101001011",
    844 => "001101001100",
    845 => "001101001101",
    846 => "001101001110",
    847 => "001101001111",
    848 => "001101010000",
    849 => "001101010001",
    850 => "001101010010",
    851 => "001101010011",
    852 => "001101010100",
    853 => "001101010101",
    854 => "001101010110",
    855 => "001101010111",
    856 => "001101011000",
    857 => "001101011001",
    858 => "001101011010",
    859 => "001101011011",
    860 => "001101011100",
    861 => "001101011101",
    862 => "001101011110",
    863 => "001101011111",
    864 => "001101100000",
    865 => "001101100001",
    866 => "001101100010",
    867 => "001101100011",
    868 => "001101100100",
    869 => "001101100101",
    870 => "001101100110",
    871 => "001101100111",
    872 => "001101101000",
    873 => "001101101001",
    874 => "001101101010",
    875 => "001101101011",
    876 => "001101101100",
    877 => "001101101101",
    878 => "001101101110",
    879 => "001101101111",
    880 => "001101110000",
    881 => "001101110001",
    882 => "001101110010",
    883 => "001101110011",
    884 => "001101110100",
    885 => "001101110101",
    886 => "001101110110",
    887 => "001101110111",
    888 => "001101111000",
    889 => "001101111001",
    890 => "001101111010",
    891 => "001101111011",
    892 => "001101111100",
    893 => "001101111101",
    894 => "001101111110",
    895 => "001101111111",
    896 => "001110000000",
    897 => "001110000001",
    898 => "001110000010",
    899 => "001110000011",
    900 => "001110000100",
    901 => "001110000101",
    902 => "001110000110",
    903 => "001110000111",
    904 => "001110001000",
    905 => "001110001001",
    906 => "001110001010",
    907 => "001110001011",
    908 => "001110001100",
    909 => "001110001101",
    910 => "001110001110",
    911 => "001110001111",
    912 => "001110010000",
    913 => "001110010001",
    914 => "001110010010",
    915 => "001110010011",
    916 => "001110010100",
    917 => "001110010101",
    918 => "001110010110",
    919 => "001110010111",
    920 => "001110011000",
    921 => "001110011001",
    922 => "001110011010",
    923 => "001110011011",
    924 => "001110011100",
    925 => "001110011101",
    926 => "001110011110",
    927 => "001110011111",
    928 => "001110100000",
    929 => "001110100001",
    930 => "001110100010",
    931 => "001110100011",
    932 => "001110100100",
    933 => "001110100101",
    934 => "001110100110",
    935 => "001110100111",
    936 => "001110101000",
    937 => "001110101001",
    938 => "001110101010",
    939 => "001110101011",
    940 => "001110101100",
    941 => "001110101101",
    942 => "001110101110",
    943 => "001110101111",
    944 => "001110110000",
    945 => "001110110001",
    946 => "001110110010",
    947 => "001110110011",
    948 => "001110110100",
    949 => "001110110101",
    950 => "001110110110",
    951 => "001110110111",
    952 => "001110111000",
    953 => "001110111001",
    954 => "001110111010",
    955 => "001110111011",
    956 => "001110111100",
    957 => "001110111101",
    958 => "001110111110",
    959 => "001110111111",
    960 => "001111000000",
    961 => "001111000001",
    962 => "001111000010",
    963 => "001111000011",
    964 => "001111000100",
    965 => "001111000101",
    966 => "001111000110",
    967 => "001111000111",
    968 => "001111001000",
    969 => "001111001001",
    970 => "001111001010",
    971 => "001111001011",
    972 => "001111001100",
    973 => "001111001101",
    974 => "001111001110",
    975 => "001111001111",
    976 => "001111010000",
    977 => "001111010001",
    978 => "001111010010",
    979 => "001111010011",
    980 => "001111010100",
    981 => "001111010101",
    982 => "001111010110",
    983 => "001111010111",
    984 => "001111011000",
    985 => "001111011001",
    986 => "001111011010",
    987 => "001111011011",
    988 => "001111011100",
    989 => "001111011101",
    990 => "001111011110",
    991 => "001111011111",
    992 => "001111100000",
    993 => "001111100001",
    994 => "001111100010",
    995 => "001111100011",
    996 => "001111100100",
    997 => "001111100101",
    998 => "001111100110",
    999 => "001111100111",
    1000 => "001111101000",
    1001 => "001111101001",
    1002 => "001111101010",
    1003 => "001111101011",
    1004 => "001111101100",
    1005 => "001111101101",
    1006 => "001111101110",
    1007 => "001111101111",
    1008 => "001111110000",
    1009 => "001111110001",
    1010 => "001111110010",
    1011 => "001111110011",
    1012 => "001111110100",
    1013 => "001111110101",
    1014 => "001111110110",
    1015 => "001111110111",
    1016 => "001111111000",
    1017 => "001111111001",
    1018 => "001111111010",
    1019 => "001111111011",
    1020 => "001111111100",
    1021 => "001111111101",
    1022 => "001111111110",
    1023 => "001111111111",
    1024 => "010000000000",
    1025 => "010000000001",
    1026 => "010000000010",
    1027 => "010000000011",
    1028 => "010000000100",
    1029 => "010000000101",
    1030 => "010000000110",
    1031 => "010000000111",
    1032 => "010000001000",
    1033 => "010000001001",
    1034 => "010000001010",
    1035 => "010000001011",
    1036 => "010000001100",
    1037 => "010000001101",
    1038 => "010000001110",
    1039 => "010000001111",
    1040 => "010000010000",
    1041 => "010000010001",
    1042 => "010000010010",
    1043 => "010000010011",
    1044 => "010000010100",
    1045 => "010000010101",
    1046 => "010000010110",
    1047 => "010000010111",
    1048 => "010000011000",
    1049 => "010000011001",
    1050 => "010000011010",
    1051 => "010000011011",
    1052 => "010000011100",
    1053 => "010000011101",
    1054 => "010000011110",
    1055 => "010000011111",
    1056 => "010000100000",
    1057 => "010000100001",
    1058 => "010000100010",
    1059 => "010000100011",
    1060 => "010000100100",
    1061 => "010000100101",
    1062 => "010000100110",
    1063 => "010000100111",
    1064 => "010000101000",
    1065 => "010000101001",
    1066 => "010000101010",
    1067 => "010000101011",
    1068 => "010000101100",
    1069 => "010000101101",
    1070 => "010000101110",
    1071 => "010000101111",
    1072 => "010000110000",
    1073 => "010000110001",
    1074 => "010000110010",
    1075 => "010000110011",
    1076 => "010000110100",
    1077 => "010000110101",
    1078 => "010000110110",
    1079 => "010000110111",
    1080 => "010000111000",
    1081 => "010000111001",
    1082 => "010000111010",
    1083 => "010000111011",
    1084 => "010000111100",
    1085 => "010000111101",
    1086 => "010000111110",
    1087 => "010000111111",
    1088 => "010001000000",
    1089 => "010001000001",
    1090 => "010001000010",
    1091 => "010001000011",
    1092 => "010001000100",
    1093 => "010001000101",
    1094 => "010001000110",
    1095 => "010001000111",
    1096 => "010001001000",
    1097 => "010001001001",
    1098 => "010001001010",
    1099 => "010001001011",
    1100 => "010001001100",
    1101 => "010001001101",
    1102 => "010001001110",
    1103 => "010001001111",
    1104 => "010001010000",
    1105 => "010001010001",
    1106 => "010001010010",
    1107 => "010001010011",
    1108 => "010001010100",
    1109 => "010001010101",
    1110 => "010001010110",
    1111 => "010001010111",
    1112 => "010001011000",
    1113 => "010001011001",
    1114 => "010001011010",
    1115 => "010001011011",
    1116 => "010001011100",
    1117 => "010001011101",
    1118 => "010001011110",
    1119 => "010001011111",
    1120 => "010001100000",
    1121 => "010001100001",
    1122 => "010001100010",
    1123 => "010001100011",
    1124 => "010001100100",
    1125 => "010001100101",
    1126 => "010001100110",
    1127 => "010001100111",
    1128 => "010001101000",
    1129 => "010001101001",
    1130 => "010001101010",
    1131 => "010001101011",
    1132 => "010001101100",
    1133 => "010001101101",
    1134 => "010001101110",
    1135 => "010001101111",
    1136 => "010001110000",
    1137 => "010001110001",
    1138 => "010001110010",
    1139 => "010001110011",
    1140 => "010001110100",
    1141 => "010001110101",
    1142 => "010001110110",
    1143 => "010001110111",
    1144 => "010001111000",
    1145 => "010001111001",
    1146 => "010001111010",
    1147 => "010001111011",
    1148 => "010001111100",
    1149 => "010001111101",
    1150 => "010001111110",
    1151 => "010001111111",
    1152 => "010010000000",
    1153 => "010010000001",
    1154 => "010010000010",
    1155 => "010010000011",
    1156 => "010010000100",
    1157 => "010010000101",
    1158 => "010010000110",
    1159 => "010010000111",
    1160 => "010010001000",
    1161 => "010010001001",
    1162 => "010010001010",
    1163 => "010010001011",
    1164 => "010010001100",
    1165 => "010010001101",
    1166 => "010010001110",
    1167 => "010010001111",
    1168 => "010010010000",
    1169 => "010010010001",
    1170 => "010010010010",
    1171 => "010010010011",
    1172 => "010010010100",
    1173 => "010010010101",
    1174 => "010010010110",
    1175 => "010010010111",
    1176 => "010010011000",
    1177 => "010010011001",
    1178 => "010010011010",
    1179 => "010010011011",
    1180 => "010010011100",
    1181 => "010010011101",
    1182 => "010010011110",
    1183 => "010010011111",
    1184 => "010010100000",
    1185 => "010010100001",
    1186 => "010010100010",
    1187 => "010010100011",
    1188 => "010010100100",
    1189 => "010010100101",
    1190 => "010010100110",
    1191 => "010010100111",
    1192 => "010010101000",
    1193 => "010010101001",
    1194 => "010010101010",
    1195 => "010010101011",
    1196 => "010010101100",
    1197 => "010010101101",
    1198 => "010010101110",
    1199 => "010010101111",
    1200 => "010010110000",
    1201 => "010010110001",
    1202 => "010010110010",
    1203 => "010010110011",
    1204 => "010010110100",
    1205 => "010010110101",
    1206 => "010010110110",
    1207 => "010010110111",
    1208 => "010010111000",
    1209 => "010010111001",
    1210 => "010010111010",
    1211 => "010010111011",
    1212 => "010010111100",
    1213 => "010010111101",
    1214 => "010010111110",
    1215 => "010010111111",
    1216 => "010011000000",
    1217 => "010011000001",
    1218 => "010011000010",
    1219 => "010011000011",
    1220 => "010011000100",
    1221 => "010011000101",
    1222 => "010011000110",
    1223 => "010011000111",
    1224 => "010011001000",
    1225 => "010011001001",
    1226 => "010011001010",
    1227 => "010011001011",
    1228 => "010011001100",
    1229 => "010011001101",
    1230 => "010011001110",
    1231 => "010011001111",
    1232 => "010011010000",
    1233 => "010011010001",
    1234 => "010011010010",
    1235 => "010011010011",
    1236 => "010011010100",
    1237 => "010011010101",
    1238 => "010011010110",
    1239 => "010011010111",
    1240 => "010011011000",
    1241 => "010011011001",
    1242 => "010011011010",
    1243 => "010011011011",
    1244 => "010011011100",
    1245 => "010011011101",
    1246 => "010011011110",
    1247 => "010011011111",
    1248 => "010011100000",
    1249 => "010011100001",
    1250 => "010011100010",
    1251 => "010011100011",
    1252 => "010011100100",
    1253 => "010011100101",
    1254 => "010011100110",
    1255 => "010011100111",
    1256 => "010011101000",
    1257 => "010011101001",
    1258 => "010011101010",
    1259 => "010011101011",
    1260 => "010011101100",
    1261 => "010011101101",
    1262 => "010011101110",
    1263 => "010011101111",
    1264 => "010011110000",
    1265 => "010011110001",
    1266 => "010011110010",
    1267 => "010011110011",
    1268 => "010011110100",
    1269 => "010011110101",
    1270 => "010011110110",
    1271 => "010011110111",
    1272 => "010011111000",
    1273 => "010011111001",
    1274 => "010011111010",
    1275 => "010011111011",
    1276 => "010011111100",
    1277 => "010011111101",
    1278 => "010011111110",
    1279 => "010011111111",
    1280 => "010100000000",
    1281 => "010100000001",
    1282 => "010100000010",
    1283 => "010100000011",
    1284 => "010100000100",
    1285 => "010100000101",
    1286 => "010100000110",
    1287 => "010100000111",
    1288 => "010100001000",
    1289 => "010100001001",
    1290 => "010100001010",
    1291 => "010100001011",
    1292 => "010100001100",
    1293 => "010100001101",
    1294 => "010100001110",
    1295 => "010100001111",
    1296 => "010100010000",
    1297 => "010100010001",
    1298 => "010100010010",
    1299 => "010100010011",
    1300 => "010100010100",
    1301 => "010100010101",
    1302 => "010100010110",
    1303 => "010100010111",
    1304 => "010100011000",
    1305 => "010100011001",
    1306 => "010100011010",
    1307 => "010100011011",
    1308 => "010100011100",
    1309 => "010100011101",
    1310 => "010100011110",
    1311 => "010100011111",
    1312 => "010100100000",
    1313 => "010100100001",
    1314 => "010100100010",
    1315 => "010100100011",
    1316 => "010100100100",
    1317 => "010100100101",
    1318 => "010100100110",
    1319 => "010100100111",
    1320 => "010100101000",
    1321 => "010100101001",
    1322 => "010100101010",
    1323 => "010100101011",
    1324 => "010100101100",
    1325 => "010100101101",
    1326 => "010100101110",
    1327 => "010100101111",
    1328 => "010100110000",
    1329 => "010100110001",
    1330 => "010100110010",
    1331 => "010100110011",
    1332 => "010100110100",
    1333 => "010100110101",
    1334 => "010100110110",
    1335 => "010100110111",
    1336 => "010100111000",
    1337 => "010100111001",
    1338 => "010100111010",
    1339 => "010100111011",
    1340 => "010100111100",
    1341 => "010100111101",
    1342 => "010100111110",
    1343 => "010100111111",
    1344 => "010101000000",
    1345 => "010101000001",
    1346 => "010101000010",
    1347 => "010101000011",
    1348 => "010101000100",
    1349 => "010101000101",
    1350 => "010101000110",
    1351 => "010101000111",
    1352 => "010101001000",
    1353 => "010101001001",
    1354 => "010101001010",
    1355 => "010101001011",
    1356 => "010101001100",
    1357 => "010101001101",
    1358 => "010101001110",
    1359 => "010101001111",
    1360 => "010101010000",
    1361 => "010101010001",
    1362 => "010101010010",
    1363 => "010101010011",
    1364 => "010101010100",
    1365 => "010101010101",
    1366 => "010101010110",
    1367 => "010101010111",
    1368 => "010101011000",
    1369 => "010101011001",
    1370 => "010101011010",
    1371 => "010101011011",
    1372 => "010101011100",
    1373 => "010101011101",
    1374 => "010101011110",
    1375 => "010101011111",
    1376 => "010101100000",
    1377 => "010101100001",
    1378 => "010101100010",
    1379 => "010101100011",
    1380 => "010101100100",
    1381 => "010101100101",
    1382 => "010101100110",
    1383 => "010101100111",
    1384 => "010101101000",
    1385 => "010101101001",
    1386 => "010101101010",
    1387 => "010101101011",
    1388 => "010101101100",
    1389 => "010101101101",
    1390 => "010101101110",
    1391 => "010101101111",
    1392 => "010101110000",
    1393 => "010101110001",
    1394 => "010101110010",
    1395 => "010101110011",
    1396 => "010101110100",
    1397 => "010101110101",
    1398 => "010101110110",
    1399 => "010101110111",
    1400 => "010101111000",
    1401 => "010101111001",
    1402 => "010101111010",
    1403 => "010101111011",
    1404 => "010101111100",
    1405 => "010101111101",
    1406 => "010101111110",
    1407 => "010101111111",
    1408 => "010110000000",
    1409 => "010110000001",
    1410 => "010110000010",
    1411 => "010110000011",
    1412 => "010110000100",
    1413 => "010110000101",
    1414 => "010110000110",
    1415 => "010110000111",
    1416 => "010110001000",
    1417 => "010110001001",
    1418 => "010110001010",
    1419 => "010110001011",
    1420 => "010110001100",
    1421 => "010110001101",
    1422 => "010110001110",
    1423 => "010110001111",
    1424 => "010110010000",
    1425 => "010110010001",
    1426 => "010110010010",
    1427 => "010110010011",
    1428 => "010110010100",
    1429 => "010110010101",
    1430 => "010110010110",
    1431 => "010110010111",
    1432 => "010110011000",
    1433 => "010110011001",
    1434 => "010110011010",
    1435 => "010110011011",
    1436 => "010110011100",
    1437 => "010110011101",
    1438 => "010110011110",
    1439 => "010110011111",
    1440 => "010110100000",
    1441 => "010110100001",
    1442 => "010110100010",
    1443 => "010110100011",
    1444 => "010110100100",
    1445 => "010110100101",
    1446 => "010110100110",
    1447 => "010110100111",
    1448 => "010110101000",
    1449 => "010110101001",
    1450 => "010110101010",
    1451 => "010110101011",
    1452 => "010110101100",
    1453 => "010110101101",
    1454 => "010110101110",
    1455 => "010110101111",
    1456 => "010110110000",
    1457 => "010110110001",
    1458 => "010110110010",
    1459 => "010110110011",
    1460 => "010110110100",
    1461 => "010110110101",
    1462 => "010110110110",
    1463 => "010110110111",
    1464 => "010110111000",
    1465 => "010110111001",
    1466 => "010110111010",
    1467 => "010110111011",
    1468 => "010110111100",
    1469 => "010110111101",
    1470 => "010110111110",
    1471 => "010110111111",
    1472 => "010111000000",
    1473 => "010111000001",
    1474 => "010111000010",
    1475 => "010111000011",
    1476 => "010111000100",
    1477 => "010111000101",
    1478 => "010111000110",
    1479 => "010111000111",
    1480 => "010111001000",
    1481 => "010111001001",
    1482 => "010111001010",
    1483 => "010111001011",
    1484 => "010111001100",
    1485 => "010111001101",
    1486 => "010111001110",
    1487 => "010111001111",
    1488 => "010111010000",
    1489 => "010111010001",
    1490 => "010111010010",
    1491 => "010111010011",
    1492 => "010111010100",
    1493 => "010111010101",
    1494 => "010111010110",
    1495 => "010111010111",
    1496 => "010111011000",
    1497 => "010111011001",
    1498 => "010111011010",
    1499 => "010111011011",
    1500 => "010111011100",
    1501 => "010111011101",
    1502 => "010111011110",
    1503 => "010111011111",
    1504 => "010111100000",
    1505 => "010111100001",
    1506 => "010111100010",
    1507 => "010111100011",
    1508 => "010111100100",
    1509 => "010111100101",
    1510 => "010111100110",
    1511 => "010111100111",
    1512 => "010111101000",
    1513 => "010111101001",
    1514 => "010111101010",
    1515 => "010111101011",
    1516 => "010111101100",
    1517 => "010111101101",
    1518 => "010111101110",
    1519 => "010111101111",
    1520 => "010111110000",
    1521 => "010111110001",
    1522 => "010111110010",
    1523 => "010111110011",
    1524 => "010111110100",
    1525 => "010111110101",
    1526 => "010111110110",
    1527 => "010111110111",
    1528 => "010111111000",
    1529 => "010111111001",
    1530 => "010111111010",
    1531 => "010111111011",
    1532 => "010111111100",
    1533 => "010111111101",
    1534 => "010111111110",
    1535 => "010111111111",
    1536 => "011000000000",
    1537 => "011000000001",
    1538 => "011000000010",
    1539 => "011000000011",
    1540 => "011000000100",
    1541 => "011000000101",
    1542 => "011000000110",
    1543 => "011000000111",
    1544 => "011000001000",
    1545 => "011000001001",
    1546 => "011000001010",
    1547 => "011000001011",
    1548 => "011000001100",
    1549 => "011000001101",
    1550 => "011000001110",
    1551 => "011000001111",
    1552 => "011000010000",
    1553 => "011000010001",
    1554 => "011000010010",
    1555 => "011000010011",
    1556 => "011000010100",
    1557 => "011000010101",
    1558 => "011000010110",
    1559 => "011000010111",
    1560 => "011000011000",
    1561 => "011000011001",
    1562 => "011000011010",
    1563 => "011000011011",
    1564 => "011000011100",
    1565 => "011000011101",
    1566 => "011000011110",
    1567 => "011000011111",
    1568 => "011000100000",
    1569 => "011000100001",
    1570 => "011000100010",
    1571 => "011000100011",
    1572 => "011000100100",
    1573 => "011000100101",
    1574 => "011000100110",
    1575 => "011000100111",
    1576 => "011000101000",
    1577 => "011000101001",
    1578 => "011000101010",
    1579 => "011000101011",
    1580 => "011000101100",
    1581 => "011000101101",
    1582 => "011000101110",
    1583 => "011000101111",
    1584 => "011000110000",
    1585 => "011000110001",
    1586 => "011000110010",
    1587 => "011000110011",
    1588 => "011000110100",
    1589 => "011000110101",
    1590 => "011000110110",
    1591 => "011000110111",
    1592 => "011000111000",
    1593 => "011000111001",
    1594 => "011000111010",
    1595 => "011000111011",
    1596 => "011000111100",
    1597 => "011000111101",
    1598 => "011000111110",
    1599 => "011000111111",
    1600 => "011001000000",
    1601 => "011001000001",
    1602 => "011001000010",
    1603 => "011001000011",
    1604 => "011001000100",
    1605 => "011001000101",
    1606 => "011001000110",
    1607 => "011001000111",
    1608 => "011001001000",
    1609 => "011001001001",
    1610 => "011001001010",
    1611 => "011001001011",
    1612 => "011001001100",
    1613 => "011001001101",
    1614 => "011001001110",
    1615 => "011001001111",
    1616 => "011001010000",
    1617 => "011001010001",
    1618 => "011001010010",
    1619 => "011001010011",
    1620 => "011001010100",
    1621 => "011001010101",
    1622 => "011001010110",
    1623 => "011001010111",
    1624 => "011001011000",
    1625 => "011001011001",
    1626 => "011001011010",
    1627 => "011001011011",
    1628 => "011001011100",
    1629 => "011001011101",
    1630 => "011001011110",
    1631 => "011001011111",
    1632 => "011001100000",
    1633 => "011001100001",
    1634 => "011001100010",
    1635 => "011001100011",
    1636 => "011001100100",
    1637 => "011001100101",
    1638 => "011001100110",
    1639 => "011001100111",
    1640 => "011001101000",
    1641 => "011001101001",
    1642 => "011001101010",
    1643 => "011001101011",
    1644 => "011001101100",
    1645 => "011001101101",
    1646 => "011001101110",
    1647 => "011001101111",
    1648 => "011001110000",
    1649 => "011001110001",
    1650 => "011001110010",
    1651 => "011001110011",
    1652 => "011001110100",
    1653 => "011001110101",
    1654 => "011001110110",
    1655 => "011001110111",
    1656 => "011001111000",
    1657 => "011001111001",
    1658 => "011001111010",
    1659 => "011001111011",
    1660 => "011001111100",
    1661 => "011001111101",
    1662 => "011001111110",
    1663 => "011001111111",
    1664 => "011010000000",
    1665 => "011010000001",
    1666 => "011010000010",
    1667 => "011010000011",
    1668 => "011010000100",
    1669 => "011010000101",
    1670 => "011010000110",
    1671 => "011010000111",
    1672 => "011010001000",
    1673 => "011010001001",
    1674 => "011010001010",
    1675 => "011010001011",
    1676 => "011010001100",
    1677 => "011010001101",
    1678 => "011010001110",
    1679 => "011010001111",
    1680 => "011010010000",
    1681 => "011010010001",
    1682 => "011010010010",
    1683 => "011010010011",
    1684 => "011010010100",
    1685 => "011010010101",
    1686 => "011010010110",
    1687 => "011010010111",
    1688 => "011010011000",
    1689 => "011010011001",
    1690 => "011010011010",
    1691 => "011010011011",
    1692 => "011010011100",
    1693 => "011010011101",
    1694 => "011010011110",
    1695 => "011010011111",
    1696 => "011010100000",
    1697 => "011010100001",
    1698 => "011010100010",
    1699 => "011010100011",
    1700 => "011010100100",
    1701 => "011010100101",
    1702 => "011010100110",
    1703 => "011010100111",
    1704 => "011010101000",
    1705 => "011010101001",
    1706 => "011010101010",
    1707 => "011010101011",
    1708 => "011010101100",
    1709 => "011010101101",
    1710 => "011010101110",
    1711 => "011010101111",
    1712 => "011010110000",
    1713 => "011010110001",
    1714 => "011010110010",
    1715 => "011010110011",
    1716 => "011010110100",
    1717 => "011010110101",
    1718 => "011010110110",
    1719 => "011010110111",
    1720 => "011010111000",
    1721 => "011010111001",
    1722 => "011010111010",
    1723 => "011010111011",
    1724 => "011010111100",
    1725 => "011010111101",
    1726 => "011010111110",
    1727 => "011010111111",
    1728 => "011011000000",
    1729 => "011011000001",
    1730 => "011011000010",
    1731 => "011011000011",
    1732 => "011011000100",
    1733 => "011011000101",
    1734 => "011011000110",
    1735 => "011011000111",
    1736 => "011011001000",
    1737 => "011011001001",
    1738 => "011011001010",
    1739 => "011011001011",
    1740 => "011011001100",
    1741 => "011011001101",
    1742 => "011011001110",
    1743 => "011011001111",
    1744 => "011011010000",
    1745 => "011011010001",
    1746 => "011011010010",
    1747 => "011011010011",
    1748 => "011011010100",
    1749 => "011011010101",
    1750 => "011011010110",
    1751 => "011011010111",
    1752 => "011011011000",
    1753 => "011011011001",
    1754 => "011011011010",
    1755 => "011011011011",
    1756 => "011011011100",
    1757 => "011011011101",
    1758 => "011011011110",
    1759 => "011011011111",
    1760 => "011011100000",
    1761 => "011011100001",
    1762 => "011011100010",
    1763 => "011011100011",
    1764 => "011011100100",
    1765 => "011011100101",
    1766 => "011011100110",
    1767 => "011011100111",
    1768 => "011011101000",
    1769 => "011011101001",
    1770 => "011011101010",
    1771 => "011011101011",
    1772 => "011011101100",
    1773 => "011011101101",
    1774 => "011011101110",
    1775 => "011011101111",
    1776 => "011011110000",
    1777 => "011011110001",
    1778 => "011011110010",
    1779 => "011011110011",
    1780 => "011011110100",
    1781 => "011011110101",
    1782 => "011011110110",
    1783 => "011011110111",
    1784 => "011011111000",
    1785 => "011011111001",
    1786 => "011011111010",
    1787 => "011011111011",
    1788 => "011011111100",
    1789 => "011011111101",
    1790 => "011011111110",
    1791 => "011011111111",
    1792 => "011100000000",
    1793 => "011100000001",
    1794 => "011100000010",
    1795 => "011100000011",
    1796 => "011100000100",
    1797 => "011100000101",
    1798 => "011100000110",
    1799 => "011100000111",
    1800 => "011100001000",
    1801 => "011100001001",
    1802 => "011100001010",
    1803 => "011100001011",
    1804 => "011100001100",
    1805 => "011100001101",
    1806 => "011100001110",
    1807 => "011100001111",
    1808 => "011100010000",
    1809 => "011100010001",
    1810 => "011100010010",
    1811 => "011100010011",
    1812 => "011100010100",
    1813 => "011100010101",
    1814 => "011100010110",
    1815 => "011100010111",
    1816 => "011100011000",
    1817 => "011100011001",
    1818 => "011100011010",
    1819 => "011100011011",
    1820 => "011100011100",
    1821 => "011100011101",
    1822 => "011100011110",
    1823 => "011100011111",
    1824 => "011100100000",
    1825 => "011100100001",
    1826 => "011100100010",
    1827 => "011100100011",
    1828 => "011100100100",
    1829 => "011100100101",
    1830 => "011100100110",
    1831 => "011100100111",
    1832 => "011100101000",
    1833 => "011100101001",
    1834 => "011100101010",
    1835 => "011100101011",
    1836 => "011100101100",
    1837 => "011100101101",
    1838 => "011100101110",
    1839 => "011100101111",
    1840 => "011100110000",
    1841 => "011100110001",
    1842 => "011100110010",
    1843 => "011100110011",
    1844 => "011100110100",
    1845 => "011100110101",
    1846 => "011100110110",
    1847 => "011100110111",
    1848 => "011100111000",
    1849 => "011100111001",
    1850 => "011100111010",
    1851 => "011100111011",
    1852 => "011100111100",
    1853 => "011100111101",
    1854 => "011100111110",
    1855 => "011100111111",
    1856 => "011101000000",
    1857 => "011101000001",
    1858 => "011101000010",
    1859 => "011101000011",
    1860 => "011101000100",
    1861 => "011101000101",
    1862 => "011101000110",
    1863 => "011101000111",
    1864 => "011101001000",
    1865 => "011101001001",
    1866 => "011101001010",
    1867 => "011101001011",
    1868 => "011101001100",
    1869 => "011101001101",
    1870 => "011101001110",
    1871 => "011101001111",
    1872 => "011101010000",
    1873 => "011101010001",
    1874 => "011101010010",
    1875 => "011101010011",
    1876 => "011101010100",
    1877 => "011101010101",
    1878 => "011101010110",
    1879 => "011101010111",
    1880 => "011101011000",
    1881 => "011101011001",
    1882 => "011101011010",
    1883 => "011101011011",
    1884 => "011101011100",
    1885 => "011101011101",
    1886 => "011101011110",
    1887 => "011101011111",
    1888 => "011101100000",
    1889 => "011101100001",
    1890 => "011101100010",
    1891 => "011101100011",
    1892 => "011101100100",
    1893 => "011101100101",
    1894 => "011101100110",
    1895 => "011101100111",
    1896 => "011101101000",
    1897 => "011101101001",
    1898 => "011101101010",
    1899 => "011101101011",
    1900 => "011101101100",
    1901 => "011101101101",
    1902 => "011101101110",
    1903 => "011101101111",
    1904 => "011101110000",
    1905 => "011101110001",
    1906 => "011101110010",
    1907 => "011101110011",
    1908 => "011101110100",
    1909 => "011101110101",
    1910 => "011101110110",
    1911 => "011101110111",
    1912 => "011101111000",
    1913 => "011101111001",
    1914 => "011101111010",
    1915 => "011101111011",
    1916 => "011101111100",
    1917 => "011101111101",
    1918 => "011101111110",
    1919 => "011101111111",
    1920 => "011110000000",
    1921 => "011110000001",
    1922 => "011110000010",
    1923 => "011110000011",
    1924 => "011110000100",
    1925 => "011110000101",
    1926 => "011110000110",
    1927 => "011110000111",
    1928 => "011110001000",
    1929 => "011110001001",
    1930 => "011110001010",
    1931 => "011110001011",
    1932 => "011110001100",
    1933 => "011110001101",
    1934 => "011110001110",
    1935 => "011110001111",
    1936 => "011110010000",
    1937 => "011110010001",
    1938 => "011110010010",
    1939 => "011110010011",
    1940 => "011110010100",
    1941 => "011110010101",
    1942 => "011110010110",
    1943 => "011110010111",
    1944 => "011110011000",
    1945 => "011110011001",
    1946 => "011110011010",
    1947 => "011110011011",
    1948 => "011110011100",
    1949 => "011110011101",
    1950 => "011110011110",
    1951 => "011110011111",
    1952 => "011110100000",
    1953 => "011110100001",
    1954 => "011110100010",
    1955 => "011110100011",
    1956 => "011110100100",
    1957 => "011110100101",
    1958 => "011110100110",
    1959 => "011110100111",
    1960 => "011110101000",
    1961 => "011110101001",
    1962 => "011110101010",
    1963 => "011110101011",
    1964 => "011110101100",
    1965 => "011110101101",
    1966 => "011110101110",
    1967 => "011110101111",
    1968 => "011110110000",
    1969 => "011110110001",
    1970 => "011110110010",
    1971 => "011110110011",
    1972 => "011110110100",
    1973 => "011110110101",
    1974 => "011110110110",
    1975 => "011110110111",
    1976 => "011110111000",
    1977 => "011110111001",
    1978 => "011110111010",
    1979 => "011110111011",
    1980 => "011110111100",
    1981 => "011110111101",
    1982 => "011110111110",
    1983 => "011110111111",
    1984 => "011111000000",
    1985 => "011111000001",
    1986 => "011111000010",
    1987 => "011111000011",
    1988 => "011111000100",
    1989 => "011111000101",
    1990 => "011111000110",
    1991 => "011111000111",
    1992 => "011111001000",
    1993 => "011111001001",
    1994 => "011111001010",
    1995 => "011111001011",
    1996 => "011111001100",
    1997 => "011111001101",
    1998 => "011111001110",
    1999 => "011111001111",
    2000 => "011111010000",
    2001 => "011111010001",
    2002 => "011111010010",
    2003 => "011111010011",
    2004 => "011111010100",
    2005 => "011111010101",
    2006 => "011111010110",
    2007 => "011111010111",
    2008 => "011111011000",
    2009 => "011111011001",
    2010 => "011111011010",
    2011 => "011111011011",
    2012 => "011111011100",
    2013 => "011111011101",
    2014 => "011111011110",
    2015 => "011111011111",
    2016 => "011111100000",
    2017 => "011111100001",
    2018 => "011111100010",
    2019 => "011111100011",
    2020 => "011111100100",
    2021 => "011111100101",
    2022 => "011111100110",
    2023 => "011111100111",
    2024 => "011111101000",
    2025 => "011111101001",
    2026 => "011111101010",
    2027 => "011111101011",
    2028 => "011111101100",
    2029 => "011111101101",
    2030 => "011111101110",
    2031 => "011111101111",
    2032 => "011111110000",
    2033 => "011111110001",
    2034 => "011111110010",
    2035 => "011111110011",
    2036 => "011111110100",
    2037 => "011111110101",
    2038 => "011111110110",
    2039 => "011111110111",
    2040 => "011111111000",
    2041 => "011111111001",
    2042 => "011111111010",
    2043 => "011111111011",
    2044 => "011111111100",
    2045 => "011111111101",
    2046 => "011111111110",
    2047 => "011111111111",
    2048 => "100000000000",
    2049 => "100000000001",
    2050 => "100000000010",
    2051 => "100000000011",
    2052 => "100000000100",
    2053 => "100000000101",
    2054 => "100000000110",
    2055 => "100000000111",
    2056 => "100000001000",
    2057 => "100000001001",
    2058 => "100000001010",
    2059 => "100000001011",
    2060 => "100000001100",
    2061 => "100000001101",
    2062 => "100000001110",
    2063 => "100000001111",
    2064 => "100000010000",
    2065 => "100000010001",
    2066 => "100000010010",
    2067 => "100000010011",
    2068 => "100000010100",
    2069 => "100000010101",
    2070 => "100000010110",
    2071 => "100000010111",
    2072 => "100000011000",
    2073 => "100000011001",
    2074 => "100000011010",
    2075 => "100000011011",
    2076 => "100000011100",
    2077 => "100000011101",
    2078 => "100000011110",
    2079 => "100000011111",
    2080 => "100000100000",
    2081 => "100000100001",
    2082 => "100000100010",
    2083 => "100000100011",
    2084 => "100000100100",
    2085 => "100000100101",
    2086 => "100000100110",
    2087 => "100000100111",
    2088 => "100000101000",
    2089 => "100000101001",
    2090 => "100000101010",
    2091 => "100000101011",
    2092 => "100000101100",
    2093 => "100000101101",
    2094 => "100000101110",
    2095 => "100000101111",
    2096 => "100000110000",
    2097 => "100000110001",
    2098 => "100000110010",
    2099 => "100000110011",
    2100 => "100000110100",
    2101 => "100000110101",
    2102 => "100000110110",
    2103 => "100000110111",
    2104 => "100000111000",
    2105 => "100000111001",
    2106 => "100000111010",
    2107 => "100000111011",
    2108 => "100000111100",
    2109 => "100000111101",
    2110 => "100000111110",
    2111 => "100000111111",
    2112 => "100001000000",
    2113 => "100001000001",
    2114 => "100001000010",
    2115 => "100001000011",
    2116 => "100001000100",
    2117 => "100001000101",
    2118 => "100001000110",
    2119 => "100001000111",
    2120 => "100001001000",
    2121 => "100001001001",
    2122 => "100001001010",
    2123 => "100001001011",
    2124 => "100001001100",
    2125 => "100001001101",
    2126 => "100001001110",
    2127 => "100001001111",
    2128 => "100001010000",
    2129 => "100001010001",
    2130 => "100001010010",
    2131 => "100001010011",
    2132 => "100001010100",
    2133 => "100001010101",
    2134 => "100001010110",
    2135 => "100001010111",
    2136 => "100001011000",
    2137 => "100001011001",
    2138 => "100001011010",
    2139 => "100001011011",
    2140 => "100001011100",
    2141 => "100001011101",
    2142 => "100001011110",
    2143 => "100001011111",
    2144 => "100001100000",
    2145 => "100001100001",
    2146 => "100001100010",
    2147 => "100001100011",
    2148 => "100001100100",
    2149 => "100001100101",
    2150 => "100001100110",
    2151 => "100001100111",
    2152 => "100001101000",
    2153 => "100001101001",
    2154 => "100001101010",
    2155 => "100001101011",
    2156 => "100001101100",
    2157 => "100001101101",
    2158 => "100001101110",
    2159 => "100001101111",
    2160 => "100001110000",
    2161 => "100001110001",
    2162 => "100001110010",
    2163 => "100001110011",
    2164 => "100001110100",
    2165 => "100001110101",
    2166 => "100001110110",
    2167 => "100001110111",
    2168 => "100001111000",
    2169 => "100001111001",
    2170 => "100001111010",
    2171 => "100001111011",
    2172 => "100001111100",
    2173 => "100001111101",
    2174 => "100001111110",
    2175 => "100001111111",
    2176 => "100010000000",
    2177 => "100010000001",
    2178 => "100010000010",
    2179 => "100010000011",
    2180 => "100010000100",
    2181 => "100010000101",
    2182 => "100010000110",
    2183 => "100010000111",
    2184 => "100010001000",
    2185 => "100010001001",
    2186 => "100010001010",
    2187 => "100010001011",
    2188 => "100010001100",
    2189 => "100010001101",
    2190 => "100010001110",
    2191 => "100010001111",
    2192 => "100010010000",
    2193 => "100010010001",
    2194 => "100010010010",
    2195 => "100010010011",
    2196 => "100010010100",
    2197 => "100010010101",
    2198 => "100010010110",
    2199 => "100010010111",
    2200 => "100010011000",
    2201 => "100010011001",
    2202 => "100010011010",
    2203 => "100010011011",
    2204 => "100010011100",
    2205 => "100010011101",
    2206 => "100010011110",
    2207 => "100010011111",
    2208 => "100010100000",
    2209 => "100010100001",
    2210 => "100010100010",
    2211 => "100010100011",
    2212 => "100010100100",
    2213 => "100010100101",
    2214 => "100010100110",
    2215 => "100010100111",
    2216 => "100010101000",
    2217 => "100010101001",
    2218 => "100010101010",
    2219 => "100010101011",
    2220 => "100010101100",
    2221 => "100010101101",
    2222 => "100010101110",
    2223 => "100010101111",
    2224 => "100010110000",
    2225 => "100010110001",
    2226 => "100010110010",
    2227 => "100010110011",
    2228 => "100010110100",
    2229 => "100010110101",
    2230 => "100010110110",
    2231 => "100010110111",
    2232 => "100010111000",
    2233 => "100010111001",
    2234 => "100010111010",
    2235 => "100010111011",
    2236 => "100010111100",
    2237 => "100010111101",
    2238 => "100010111110",
    2239 => "100010111111",
    2240 => "100011000000",
    2241 => "100011000001",
    2242 => "100011000010",
    2243 => "100011000011",
    2244 => "100011000100",
    2245 => "100011000101",
    2246 => "100011000110",
    2247 => "100011000111",
    2248 => "100011001000",
    2249 => "100011001001",
    2250 => "100011001010",
    2251 => "100011001011",
    2252 => "100011001100",
    2253 => "100011001101",
    2254 => "100011001110",
    2255 => "100011001111",
    2256 => "100011010000",
    2257 => "100011010001",
    2258 => "100011010010",
    2259 => "100011010011",
    2260 => "100011010100",
    2261 => "100011010101",
    2262 => "100011010110",
    2263 => "100011010111",
    2264 => "100011011000",
    2265 => "100011011001",
    2266 => "100011011010",
    2267 => "100011011011",
    2268 => "100011011100",
    2269 => "100011011101",
    2270 => "100011011110",
    2271 => "100011011111",
    2272 => "100011100000",
    2273 => "100011100001",
    2274 => "100011100010",
    2275 => "100011100011",
    2276 => "100011100100",
    2277 => "100011100101",
    2278 => "100011100110",
    2279 => "100011100111",
    2280 => "100011101000",
    2281 => "100011101001",
    2282 => "100011101010",
    2283 => "100011101011",
    2284 => "100011101100",
    2285 => "100011101101",
    2286 => "100011101110",
    2287 => "100011101111",
    2288 => "100011110000",
    2289 => "100011110001",
    2290 => "100011110010",
    2291 => "100011110011",
    2292 => "100011110100",
    2293 => "100011110101",
    2294 => "100011110110",
    2295 => "100011110111",
    2296 => "100011111000",
    2297 => "100011111001",
    2298 => "100011111010",
    2299 => "100011111011",
    2300 => "100011111100",
    2301 => "100011111101",
    2302 => "100011111110",
    2303 => "100011111111",
    2304 => "100100000000",
    2305 => "100100000001",
    2306 => "100100000010",
    2307 => "100100000011",
    2308 => "100100000100",
    2309 => "100100000101",
    2310 => "100100000110",
    2311 => "100100000111",
    2312 => "100100001000",
    2313 => "100100001001",
    2314 => "100100001010",
    2315 => "100100001011",
    2316 => "100100001100",
    2317 => "100100001101",
    2318 => "100100001110",
    2319 => "100100001111",
    2320 => "100100010000",
    2321 => "100100010001",
    2322 => "100100010010",
    2323 => "100100010011",
    2324 => "100100010100",
    2325 => "100100010101",
    2326 => "100100010110",
    2327 => "100100010111",
    2328 => "100100011000",
    2329 => "100100011001",
    2330 => "100100011010",
    2331 => "100100011011",
    2332 => "100100011100",
    2333 => "100100011101",
    2334 => "100100011110",
    2335 => "100100011111",
    2336 => "100100100000",
    2337 => "100100100001",
    2338 => "100100100010",
    2339 => "100100100011",
    2340 => "100100100100",
    2341 => "100100100101",
    2342 => "100100100110",
    2343 => "100100100111",
    2344 => "100100101000",
    2345 => "100100101001",
    2346 => "100100101010",
    2347 => "100100101011",
    2348 => "100100101100",
    2349 => "100100101101",
    2350 => "100100101110",
    2351 => "100100101111",
    2352 => "100100110000",
    2353 => "100100110001",
    2354 => "100100110010",
    2355 => "100100110011",
    2356 => "100100110100",
    2357 => "100100110101",
    2358 => "100100110110",
    2359 => "100100110111",
    2360 => "100100111000",
    2361 => "100100111001",
    2362 => "100100111010",
    2363 => "100100111011",
    2364 => "100100111100",
    2365 => "100100111101",
    2366 => "100100111110",
    2367 => "100100111111",
    2368 => "100101000000",
    2369 => "100101000001",
    2370 => "100101000010",
    2371 => "100101000011",
    2372 => "100101000100",
    2373 => "100101000101",
    2374 => "100101000110",
    2375 => "100101000111",
    2376 => "100101001000",
    2377 => "100101001001",
    2378 => "100101001010",
    2379 => "100101001011",
    2380 => "100101001100",
    2381 => "100101001101",
    2382 => "100101001110",
    2383 => "100101001111",
    2384 => "100101010000",
    2385 => "100101010001",
    2386 => "100101010010",
    2387 => "100101010011",
    2388 => "100101010100",
    2389 => "100101010101",
    2390 => "100101010110",
    2391 => "100101010111",
    2392 => "100101011000",
    2393 => "100101011001",
    2394 => "100101011010",
    2395 => "100101011011",
    2396 => "100101011100",
    2397 => "100101011101",
    2398 => "100101011110",
    2399 => "100101011111",
    2400 => "100101100000",
    2401 => "100101100001",
    2402 => "100101100010",
    2403 => "100101100011",
    2404 => "100101100100",
    2405 => "100101100101",
    2406 => "100101100110",
    2407 => "100101100111",
    2408 => "100101101000",
    2409 => "100101101001",
    2410 => "100101101010",
    2411 => "100101101011",
    2412 => "100101101100",
    2413 => "100101101101",
    2414 => "100101101110",
    2415 => "100101101111",
    2416 => "100101110000",
    2417 => "100101110001",
    2418 => "100101110010",
    2419 => "100101110011",
    2420 => "100101110100",
    2421 => "100101110101",
    2422 => "100101110110",
    2423 => "100101110111",
    2424 => "100101111000",
    2425 => "100101111001",
    2426 => "100101111010",
    2427 => "100101111011",
    2428 => "100101111100",
    2429 => "100101111101",
    2430 => "100101111110",
    2431 => "100101111111",
    2432 => "100110000000",
    2433 => "100110000001",
    2434 => "100110000010",
    2435 => "100110000011",
    2436 => "100110000100",
    2437 => "100110000101",
    2438 => "100110000110",
    2439 => "100110000111",
    2440 => "100110001000",
    2441 => "100110001001",
    2442 => "100110001010",
    2443 => "100110001011",
    2444 => "100110001100",
    2445 => "100110001101",
    2446 => "100110001110",
    2447 => "100110001111",
    2448 => "100110010000",
    2449 => "100110010001",
    2450 => "100110010010",
    2451 => "100110010011",
    2452 => "100110010100",
    2453 => "100110010101",
    2454 => "100110010110",
    2455 => "100110010111",
    2456 => "100110011000",
    2457 => "100110011001",
    2458 => "100110011010",
    2459 => "100110011011",
    2460 => "100110011100",
    2461 => "100110011101",
    2462 => "100110011110",
    2463 => "100110011111",
    2464 => "100110100000",
    2465 => "100110100001",
    2466 => "100110100010",
    2467 => "100110100011",
    2468 => "100110100100",
    2469 => "100110100101",
    2470 => "100110100110",
    2471 => "100110100111",
    2472 => "100110101000",
    2473 => "100110101001",
    2474 => "100110101010",
    2475 => "100110101011",
    2476 => "100110101100",
    2477 => "100110101101",
    2478 => "100110101110",
    2479 => "100110101111",
    2480 => "100110110000",
    2481 => "100110110001",
    2482 => "100110110010",
    2483 => "100110110011",
    2484 => "100110110100",
    2485 => "100110110101",
    2486 => "100110110110",
    2487 => "100110110111",
    2488 => "100110111000",
    2489 => "100110111001",
    2490 => "100110111010",
    2491 => "100110111011",
    2492 => "100110111100",
    2493 => "100110111101",
    2494 => "100110111110",
    2495 => "100110111111",
    2496 => "100111000000",
    2497 => "100111000001",
    2498 => "100111000010",
    2499 => "100111000011",
    2500 => "100111000100",
    2501 => "100111000101",
    2502 => "100111000110",
    2503 => "100111000111",
    2504 => "100111001000",
    2505 => "100111001001",
    2506 => "100111001010",
    2507 => "100111001011",
    2508 => "100111001100",
    2509 => "100111001101",
    2510 => "100111001110",
    2511 => "100111001111",
    2512 => "100111010000",
    2513 => "100111010001",
    2514 => "100111010010",
    2515 => "100111010011",
    2516 => "100111010100",
    2517 => "100111010101",
    2518 => "100111010110",
    2519 => "100111010111",
    2520 => "100111011000",
    2521 => "100111011001",
    2522 => "100111011010",
    2523 => "100111011011",
    2524 => "100111011100",
    2525 => "100111011101",
    2526 => "100111011110",
    2527 => "100111011111",
    2528 => "100111100000",
    2529 => "100111100001",
    2530 => "100111100010",
    2531 => "100111100011",
    2532 => "100111100100",
    2533 => "100111100101",
    2534 => "100111100110",
    2535 => "100111100111",
    2536 => "100111101000",
    2537 => "100111101001",
    2538 => "100111101010",
    2539 => "100111101011",
    2540 => "100111101100",
    2541 => "100111101101",
    2542 => "100111101110",
    2543 => "100111101111",
    2544 => "100111110000",
    2545 => "100111110001",
    2546 => "100111110010",
    2547 => "100111110011",
    2548 => "100111110100",
    2549 => "100111110101",
    2550 => "100111110110",
    2551 => "100111110111",
    2552 => "100111111000",
    2553 => "100111111001",
    2554 => "100111111010",
    2555 => "100111111011",
    2556 => "100111111100",
    2557 => "100111111101",
    2558 => "100111111110",
    2559 => "100111111111",
    2560 => "101000000000",
    2561 => "101000000001",
    2562 => "101000000010",
    2563 => "101000000011",
    2564 => "101000000100",
    2565 => "101000000101",
    2566 => "101000000110",
    2567 => "101000000111",
    2568 => "101000001000",
    2569 => "101000001001",
    2570 => "101000001010",
    2571 => "101000001011",
    2572 => "101000001100",
    2573 => "101000001101",
    2574 => "101000001110",
    2575 => "101000001111",
    2576 => "101000010000",
    2577 => "101000010001",
    2578 => "101000010010",
    2579 => "101000010011",
    2580 => "101000010100",
    2581 => "101000010101",
    2582 => "101000010110",
    2583 => "101000010111",
    2584 => "101000011000",
    2585 => "101000011001",
    2586 => "101000011010",
    2587 => "101000011011",
    2588 => "101000011100",
    2589 => "101000011101",
    2590 => "101000011110",
    2591 => "101000011111",
    2592 => "101000100000",
    2593 => "101000100001",
    2594 => "101000100010",
    2595 => "101000100011",
    2596 => "101000100100",
    2597 => "101000100101",
    2598 => "101000100110",
    2599 => "101000100111",
    2600 => "101000101000",
    2601 => "101000101001",
    2602 => "101000101010",
    2603 => "101000101011",
    2604 => "101000101100",
    2605 => "101000101101",
    2606 => "101000101110",
    2607 => "101000101111",
    2608 => "101000110000",
    2609 => "101000110001",
    2610 => "101000110010",
    2611 => "101000110011",
    2612 => "101000110100",
    2613 => "101000110101",
    2614 => "101000110110",
    2615 => "101000110111",
    2616 => "101000111000",
    2617 => "101000111001",
    2618 => "101000111010",
    2619 => "101000111011",
    2620 => "101000111100",
    2621 => "101000111101",
    2622 => "101000111110",
    2623 => "101000111111",
    2624 => "101001000000",
    2625 => "101001000001",
    2626 => "101001000010",
    2627 => "101001000011",
    2628 => "101001000100",
    2629 => "101001000101",
    2630 => "101001000110",
    2631 => "101001000111",
    2632 => "101001001000",
    2633 => "101001001001",
    2634 => "101001001010",
    2635 => "101001001011",
    2636 => "101001001100",
    2637 => "101001001101",
    2638 => "101001001110",
    2639 => "101001001111",
    2640 => "101001010000",
    2641 => "101001010001",
    2642 => "101001010010",
    2643 => "101001010011",
    2644 => "101001010100",
    2645 => "101001010101",
    2646 => "101001010110",
    2647 => "101001010111",
    2648 => "101001011000",
    2649 => "101001011001",
    2650 => "101001011010",
    2651 => "101001011011",
    2652 => "101001011100",
    2653 => "101001011101",
    2654 => "101001011110",
    2655 => "101001011111",
    2656 => "101001100000",
    2657 => "101001100001",
    2658 => "101001100010",
    2659 => "101001100011",
    2660 => "101001100100",
    2661 => "101001100101",
    2662 => "101001100110",
    2663 => "101001100111",
    2664 => "101001101000",
    2665 => "101001101001",
    2666 => "101001101010",
    2667 => "101001101011",
    2668 => "101001101100",
    2669 => "101001101101",
    2670 => "101001101110",
    2671 => "101001101111",
    2672 => "101001110000",
    2673 => "101001110001",
    2674 => "101001110010",
    2675 => "101001110011",
    2676 => "101001110100",
    2677 => "101001110101",
    2678 => "101001110110",
    2679 => "101001110111",
    2680 => "101001111000",
    2681 => "101001111001",
    2682 => "101001111010",
    2683 => "101001111011",
    2684 => "101001111100",
    2685 => "101001111101",
    2686 => "101001111110",
    2687 => "101001111111",
    2688 => "101010000000",
    2689 => "101010000001",
    2690 => "101010000010",
    2691 => "101010000011",
    2692 => "101010000100",
    2693 => "101010000101",
    2694 => "101010000110",
    2695 => "101010000111",
    2696 => "101010001000",
    2697 => "101010001001",
    2698 => "101010001010",
    2699 => "101010001011",
    2700 => "101010001100",
    2701 => "101010001101",
    2702 => "101010001110",
    2703 => "101010001111",
    2704 => "101010010000",
    2705 => "101010010001",
    2706 => "101010010010",
    2707 => "101010010011",
    2708 => "101010010100",
    2709 => "101010010101",
    2710 => "101010010110",
    2711 => "101010010111",
    2712 => "101010011000",
    2713 => "101010011001",
    2714 => "101010011010",
    2715 => "101010011011",
    2716 => "101010011100",
    2717 => "101010011101",
    2718 => "101010011110",
    2719 => "101010011111",
    2720 => "101010100000",
    2721 => "101010100001",
    2722 => "101010100010",
    2723 => "101010100011",
    2724 => "101010100100",
    2725 => "101010100101",
    2726 => "101010100110",
    2727 => "101010100111",
    2728 => "101010101000",
    2729 => "101010101001",
    2730 => "101010101010",
    2731 => "101010101011",
    2732 => "101010101100",
    2733 => "101010101101",
    2734 => "101010101110",
    2735 => "101010101111",
    2736 => "101010110000",
    2737 => "101010110001",
    2738 => "101010110010",
    2739 => "101010110011",
    2740 => "101010110100",
    2741 => "101010110101",
    2742 => "101010110110",
    2743 => "101010110111",
    2744 => "101010111000",
    2745 => "101010111001",
    2746 => "101010111010",
    2747 => "101010111011",
    2748 => "101010111100",
    2749 => "101010111101",
    2750 => "101010111110",
    2751 => "101010111111",
    2752 => "101011000000",
    2753 => "101011000001",
    2754 => "101011000010",
    2755 => "101011000011",
    2756 => "101011000100",
    2757 => "101011000101",
    2758 => "101011000110",
    2759 => "101011000111",
    2760 => "101011001000",
    2761 => "101011001001",
    2762 => "101011001010",
    2763 => "101011001011",
    2764 => "101011001100",
    2765 => "101011001101",
    2766 => "101011001110",
    2767 => "101011001111",
    2768 => "101011010000",
    2769 => "101011010001",
    2770 => "101011010010",
    2771 => "101011010011",
    2772 => "101011010100",
    2773 => "101011010101",
    2774 => "101011010110",
    2775 => "101011010111",
    2776 => "101011011000",
    2777 => "101011011001",
    2778 => "101011011010",
    2779 => "101011011011",
    2780 => "101011011100",
    2781 => "101011011101",
    2782 => "101011011110",
    2783 => "101011011111",
    2784 => "101011100000",
    2785 => "101011100001",
    2786 => "101011100010",
    2787 => "101011100011",
    2788 => "101011100100",
    2789 => "101011100101",
    2790 => "101011100110",
    2791 => "101011100111",
    2792 => "101011101000",
    2793 => "101011101001",
    2794 => "101011101010",
    2795 => "101011101011",
    2796 => "101011101100",
    2797 => "101011101101",
    2798 => "101011101110",
    2799 => "101011101111",
    2800 => "101011110000",
    2801 => "101011110001",
    2802 => "101011110010",
    2803 => "101011110011",
    2804 => "101011110100",
    2805 => "101011110101",
    2806 => "101011110110",
    2807 => "101011110111",
    2808 => "101011111000",
    2809 => "101011111001",
    2810 => "101011111010",
    2811 => "101011111011",
    2812 => "101011111100",
    2813 => "101011111101",
    2814 => "101011111110",
    2815 => "101011111111",
    2816 => "101100000000",
    2817 => "101100000001",
    2818 => "101100000010",
    2819 => "101100000011",
    2820 => "101100000100",
    2821 => "101100000101",
    2822 => "101100000110",
    2823 => "101100000111",
    2824 => "101100001000",
    2825 => "101100001001",
    2826 => "101100001010",
    2827 => "101100001011",
    2828 => "101100001100",
    2829 => "101100001101",
    2830 => "101100001110",
    2831 => "101100001111",
    2832 => "101100010000",
    2833 => "101100010001",
    2834 => "101100010010",
    2835 => "101100010011",
    2836 => "101100010100",
    2837 => "101100010101",
    2838 => "101100010110",
    2839 => "101100010111",
    2840 => "101100011000",
    2841 => "101100011001",
    2842 => "101100011010",
    2843 => "101100011011",
    2844 => "101100011100",
    2845 => "101100011101",
    2846 => "101100011110",
    2847 => "101100011111",
    2848 => "101100100000",
    2849 => "101100100001",
    2850 => "101100100010",
    2851 => "101100100011",
    2852 => "101100100100",
    2853 => "101100100101",
    2854 => "101100100110",
    2855 => "101100100111",
    2856 => "101100101000",
    2857 => "101100101001",
    2858 => "101100101010",
    2859 => "101100101011",
    2860 => "101100101100",
    2861 => "101100101101",
    2862 => "101100101110",
    2863 => "101100101111",
    2864 => "101100110000",
    2865 => "101100110001",
    2866 => "101100110010",
    2867 => "101100110011",
    2868 => "101100110100",
    2869 => "101100110101",
    2870 => "101100110110",
    2871 => "101100110111",
    2872 => "101100111000",
    2873 => "101100111001",
    2874 => "101100111010",
    2875 => "101100111011",
    2876 => "101100111100",
    2877 => "101100111101",
    2878 => "101100111110",
    2879 => "101100111111",
    2880 => "101101000000",
    2881 => "101101000001",
    2882 => "101101000010",
    2883 => "101101000011",
    2884 => "101101000100",
    2885 => "101101000101",
    2886 => "101101000110",
    2887 => "101101000111",
    2888 => "101101001000",
    2889 => "101101001001",
    2890 => "101101001010",
    2891 => "101101001011",
    2892 => "101101001100",
    2893 => "101101001101",
    2894 => "101101001110",
    2895 => "101101001111",
    2896 => "101101010000",
    2897 => "101101010001",
    2898 => "101101010010",
    2899 => "101101010011",
    2900 => "101101010100",
    2901 => "101101010101",
    2902 => "101101010110",
    2903 => "101101010111",
    2904 => "101101011000",
    2905 => "101101011001",
    2906 => "101101011010",
    2907 => "101101011011",
    2908 => "101101011100",
    2909 => "101101011101",
    2910 => "101101011110",
    2911 => "101101011111",
    2912 => "101101100000",
    2913 => "101101100001",
    2914 => "101101100010",
    2915 => "101101100011",
    2916 => "101101100100",
    2917 => "101101100101",
    2918 => "101101100110",
    2919 => "101101100111",
    2920 => "101101101000",
    2921 => "101101101001",
    2922 => "101101101010",
    2923 => "101101101011",
    2924 => "101101101100",
    2925 => "101101101101",
    2926 => "101101101110",
    2927 => "101101101111",
    2928 => "101101110000",
    2929 => "101101110001",
    2930 => "101101110010",
    2931 => "101101110011",
    2932 => "101101110100",
    2933 => "101101110101",
    2934 => "101101110110",
    2935 => "101101110111",
    2936 => "101101111000",
    2937 => "101101111001",
    2938 => "101101111010",
    2939 => "101101111011",
    2940 => "101101111100",
    2941 => "101101111101",
    2942 => "101101111110",
    2943 => "101101111111",
    2944 => "101110000000",
    2945 => "101110000001",
    2946 => "101110000010",
    2947 => "101110000011",
    2948 => "101110000100",
    2949 => "101110000101",
    2950 => "101110000110",
    2951 => "101110000111",
    2952 => "101110001000",
    2953 => "101110001001",
    2954 => "101110001010",
    2955 => "101110001011",
    2956 => "101110001100",
    2957 => "101110001101",
    2958 => "101110001110",
    2959 => "101110001111",
    2960 => "101110010000",
    2961 => "101110010001",
    2962 => "101110010010",
    2963 => "101110010011",
    2964 => "101110010100",
    2965 => "101110010101",
    2966 => "101110010110",
    2967 => "101110010111",
    2968 => "101110011000",
    2969 => "101110011001",
    2970 => "101110011010",
    2971 => "101110011011",
    2972 => "101110011100",
    2973 => "101110011101",
    2974 => "101110011110",
    2975 => "101110011111",
    2976 => "101110100000",
    2977 => "101110100001",
    2978 => "101110100010",
    2979 => "101110100011",
    2980 => "101110100100",
    2981 => "101110100101",
    2982 => "101110100110",
    2983 => "101110100111",
    2984 => "101110101000",
    2985 => "101110101001",
    2986 => "101110101010",
    2987 => "101110101011",
    2988 => "101110101100",
    2989 => "101110101101",
    2990 => "101110101110",
    2991 => "101110101111",
    2992 => "101110110000",
    2993 => "101110110001",
    2994 => "101110110010",
    2995 => "101110110011",
    2996 => "101110110100",
    2997 => "101110110101",
    2998 => "101110110110",
    2999 => "101110110111",
    3000 => "101110111000",
    3001 => "101110111001",
    3002 => "101110111010",
    3003 => "101110111011",
    3004 => "101110111100",
    3005 => "101110111101",
    3006 => "101110111110",
    3007 => "101110111111",
    3008 => "101111000000",
    3009 => "101111000001",
    3010 => "101111000010",
    3011 => "101111000011",
    3012 => "101111000100",
    3013 => "101111000101",
    3014 => "101111000110",
    3015 => "101111000111",
    3016 => "101111001000",
    3017 => "101111001001",
    3018 => "101111001010",
    3019 => "101111001011",
    3020 => "101111001100",
    3021 => "101111001101",
    3022 => "101111001110",
    3023 => "101111001111",
    3024 => "101111010000",
    3025 => "101111010001",
    3026 => "101111010010",
    3027 => "101111010011",
    3028 => "101111010100",
    3029 => "101111010101",
    3030 => "101111010110",
    3031 => "101111010111",
    3032 => "101111011000",
    3033 => "101111011001",
    3034 => "101111011010",
    3035 => "101111011011",
    3036 => "101111011100",
    3037 => "101111011101",
    3038 => "101111011110",
    3039 => "101111011111",
    3040 => "101111100000",
    3041 => "101111100001",
    3042 => "101111100010",
    3043 => "101111100011",
    3044 => "101111100100",
    3045 => "101111100101",
    3046 => "101111100110",
    3047 => "101111100111",
    3048 => "101111101000",
    3049 => "101111101001",
    3050 => "101111101010",
    3051 => "101111101011",
    3052 => "101111101100",
    3053 => "101111101101",
    3054 => "101111101110",
    3055 => "101111101111",
    3056 => "101111110000",
    3057 => "101111110001",
    3058 => "101111110010",
    3059 => "101111110011",
    3060 => "101111110100",
    3061 => "101111110101",
    3062 => "101111110110",
    3063 => "101111110111",
    3064 => "101111111000",
    3065 => "101111111001",
    3066 => "101111111010",
    3067 => "101111111011",
    3068 => "101111111100",
    3069 => "101111111101",
    3070 => "101111111110",
    3071 => "101111111111",
    3072 => "110000000000",
    3073 => "110000000001",
    3074 => "110000000010",
    3075 => "110000000011",
    3076 => "110000000100",
    3077 => "110000000101",
    3078 => "110000000110",
    3079 => "110000000111",
    3080 => "110000001000",
    3081 => "110000001001",
    3082 => "110000001010",
    3083 => "110000001011",
    3084 => "110000001100",
    3085 => "110000001101",
    3086 => "110000001110",
    3087 => "110000001111",
    3088 => "110000010000",
    3089 => "110000010001",
    3090 => "110000010010",
    3091 => "110000010011",
    3092 => "110000010100",
    3093 => "110000010101",
    3094 => "110000010110",
    3095 => "110000010111",
    3096 => "110000011000",
    3097 => "110000011001",
    3098 => "110000011010",
    3099 => "110000011011",
    3100 => "110000011100",
    3101 => "110000011101",
    3102 => "110000011110",
    3103 => "110000011111",
    3104 => "110000100000",
    3105 => "110000100001",
    3106 => "110000100010",
    3107 => "110000100011",
    3108 => "110000100100",
    3109 => "110000100101",
    3110 => "110000100110",
    3111 => "110000100111",
    3112 => "110000101000",
    3113 => "110000101001",
    3114 => "110000101010",
    3115 => "110000101011",
    3116 => "110000101100",
    3117 => "110000101101",
    3118 => "110000101110",
    3119 => "110000101111",
    3120 => "110000110000",
    3121 => "110000110001",
    3122 => "110000110010",
    3123 => "110000110011",
    3124 => "110000110100",
    3125 => "110000110101",
    3126 => "110000110110",
    3127 => "110000110111",
    3128 => "110000111000",
    3129 => "110000111001",
    3130 => "110000111010",
    3131 => "110000111011",
    3132 => "110000111100",
    3133 => "110000111101",
    3134 => "110000111110",
    3135 => "110000111111",
    3136 => "110001000000",
    3137 => "110001000001",
    3138 => "110001000010",
    3139 => "110001000011",
    3140 => "110001000100",
    3141 => "110001000101",
    3142 => "110001000110",
    3143 => "110001000111",
    3144 => "110001001000",
    3145 => "110001001001",
    3146 => "110001001010",
    3147 => "110001001011",
    3148 => "110001001100",
    3149 => "110001001101",
    3150 => "110001001110",
    3151 => "110001001111",
    3152 => "110001010000",
    3153 => "110001010001",
    3154 => "110001010010",
    3155 => "110001010011",
    3156 => "110001010100",
    3157 => "110001010101",
    3158 => "110001010110",
    3159 => "110001010111",
    3160 => "110001011000",
    3161 => "110001011001",
    3162 => "110001011010",
    3163 => "110001011011",
    3164 => "110001011100",
    3165 => "110001011101",
    3166 => "110001011110",
    3167 => "110001011111",
    3168 => "110001100000",
    3169 => "110001100001",
    3170 => "110001100010",
    3171 => "110001100011",
    3172 => "110001100100",
    3173 => "110001100101",
    3174 => "110001100110",
    3175 => "110001100111",
    3176 => "110001101000",
    3177 => "110001101001",
    3178 => "110001101010",
    3179 => "110001101011",
    3180 => "110001101100",
    3181 => "110001101101",
    3182 => "110001101110",
    3183 => "110001101111",
    3184 => "110001110000",
    3185 => "110001110001",
    3186 => "110001110010",
    3187 => "110001110011",
    3188 => "110001110100",
    3189 => "110001110101",
    3190 => "110001110110",
    3191 => "110001110111",
    3192 => "110001111000",
    3193 => "110001111001",
    3194 => "110001111010",
    3195 => "110001111011",
    3196 => "110001111100",
    3197 => "110001111101",
    3198 => "110001111110",
    3199 => "110001111111",
    3200 => "110010000000",
    3201 => "110010000001",
    3202 => "110010000010",
    3203 => "110010000011",
    3204 => "110010000100",
    3205 => "110010000101",
    3206 => "110010000110",
    3207 => "110010000111",
    3208 => "110010001000",
    3209 => "110010001001",
    3210 => "110010001010",
    3211 => "110010001011",
    3212 => "110010001100",
    3213 => "110010001101",
    3214 => "110010001110",
    3215 => "110010001111",
    3216 => "110010010000",
    3217 => "110010010001",
    3218 => "110010010010",
    3219 => "110010010011",
    3220 => "110010010100",
    3221 => "110010010101",
    3222 => "110010010110",
    3223 => "110010010111",
    3224 => "110010011000",
    3225 => "110010011001",
    3226 => "110010011010",
    3227 => "110010011011",
    3228 => "110010011100",
    3229 => "110010011101",
    3230 => "110010011110",
    3231 => "110010011111",
    3232 => "110010100000",
    3233 => "110010100001",
    3234 => "110010100010",
    3235 => "110010100011",
    3236 => "110010100100",
    3237 => "110010100101",
    3238 => "110010100110",
    3239 => "110010100111",
    3240 => "110010101000",
    3241 => "110010101001",
    3242 => "110010101010",
    3243 => "110010101011",
    3244 => "110010101100",
    3245 => "110010101101",
    3246 => "110010101110",
    3247 => "110010101111",
    3248 => "110010110000",
    3249 => "110010110001",
    3250 => "110010110010",
    3251 => "110010110011",
    3252 => "110010110100",
    3253 => "110010110101",
    3254 => "110010110110",
    3255 => "110010110111",
    3256 => "110010111000",
    3257 => "110010111001",
    3258 => "110010111010",
    3259 => "110010111011",
    3260 => "110010111100",
    3261 => "110010111101",
    3262 => "110010111110",
    3263 => "110010111111",
    3264 => "110011000000",
    3265 => "110011000001",
    3266 => "110011000010",
    3267 => "110011000011",
    3268 => "110011000100",
    3269 => "110011000101",
    3270 => "110011000110",
    3271 => "110011000111",
    3272 => "110011001000",
    3273 => "110011001001",
    3274 => "110011001010",
    3275 => "110011001011",
    3276 => "110011001100",
    3277 => "110011001101",
    3278 => "110011001110",
    3279 => "110011001111",
    3280 => "110011010000",
    3281 => "110011010001",
    3282 => "110011010010",
    3283 => "110011010011",
    3284 => "110011010100",
    3285 => "110011010101",
    3286 => "110011010110",
    3287 => "110011010111",
    3288 => "110011011000",
    3289 => "110011011001",
    3290 => "110011011010",
    3291 => "110011011011",
    3292 => "110011011100",
    3293 => "110011011101",
    3294 => "110011011110",
    3295 => "110011011111",
    3296 => "110011100000",
    3297 => "110011100001",
    3298 => "110011100010",
    3299 => "110011100011",
    3300 => "110011100100",
    3301 => "110011100101",
    3302 => "110011100110",
    3303 => "110011100111",
    3304 => "110011101000",
    3305 => "110011101001",
    3306 => "110011101010",
    3307 => "110011101011",
    3308 => "110011101100",
    3309 => "110011101101",
    3310 => "110011101110",
    3311 => "110011101111",
    3312 => "110011110000",
    3313 => "110011110001",
    3314 => "110011110010",
    3315 => "110011110011",
    3316 => "110011110100",
    3317 => "110011110101",
    3318 => "110011110110",
    3319 => "110011110111",
    3320 => "110011111000",
    3321 => "110011111001",
    3322 => "110011111010",
    3323 => "110011111011",
    3324 => "110011111100",
    3325 => "110011111101",
    3326 => "110011111110",
    3327 => "110011111111",
    3328 => "110100000000",
    3329 => "110100000001",
    3330 => "110100000010",
    3331 => "110100000011",
    3332 => "110100000100",
    3333 => "110100000101",
    3334 => "110100000110",
    3335 => "110100000111",
    3336 => "110100001000",
    3337 => "110100001001",
    3338 => "110100001010",
    3339 => "110100001011",
    3340 => "110100001100",
    3341 => "110100001101",
    3342 => "110100001110",
    3343 => "110100001111",
    3344 => "110100010000",
    3345 => "110100010001",
    3346 => "110100010010",
    3347 => "110100010011",
    3348 => "110100010100",
    3349 => "110100010101",
    3350 => "110100010110",
    3351 => "110100010111",
    3352 => "110100011000",
    3353 => "110100011001",
    3354 => "110100011010",
    3355 => "110100011011",
    3356 => "110100011100",
    3357 => "110100011101",
    3358 => "110100011110",
    3359 => "110100011111",
    3360 => "110100100000",
    3361 => "110100100001",
    3362 => "110100100010",
    3363 => "110100100011",
    3364 => "110100100100",
    3365 => "110100100101",
    3366 => "110100100110",
    3367 => "110100100111",
    3368 => "110100101000",
    3369 => "110100101001",
    3370 => "110100101010",
    3371 => "110100101011",
    3372 => "110100101100",
    3373 => "110100101101",
    3374 => "110100101110",
    3375 => "110100101111",
    3376 => "110100110000",
    3377 => "110100110001",
    3378 => "110100110010",
    3379 => "110100110011",
    3380 => "110100110100",
    3381 => "110100110101",
    3382 => "110100110110",
    3383 => "110100110111",
    3384 => "110100111000",
    3385 => "110100111001",
    3386 => "110100111010",
    3387 => "110100111011",
    3388 => "110100111100",
    3389 => "110100111101",
    3390 => "110100111110",
    3391 => "110100111111",
    3392 => "110101000000",
    3393 => "110101000001",
    3394 => "110101000010",
    3395 => "110101000011",
    3396 => "110101000100",
    3397 => "110101000101",
    3398 => "110101000110",
    3399 => "110101000111",
    3400 => "110101001000",
    3401 => "110101001001",
    3402 => "110101001010",
    3403 => "110101001011",
    3404 => "110101001100",
    3405 => "110101001101",
    3406 => "110101001110",
    3407 => "110101001111",
    3408 => "110101010000",
    3409 => "110101010001",
    3410 => "110101010010",
    3411 => "110101010011",
    3412 => "110101010100",
    3413 => "110101010101",
    3414 => "110101010110",
    3415 => "110101010111",
    3416 => "110101011000",
    3417 => "110101011001",
    3418 => "110101011010",
    3419 => "110101011011",
    3420 => "110101011100",
    3421 => "110101011101",
    3422 => "110101011110",
    3423 => "110101011111",
    3424 => "110101100000",
    3425 => "110101100001",
    3426 => "110101100010",
    3427 => "110101100011",
    3428 => "110101100100",
    3429 => "110101100101",
    3430 => "110101100110",
    3431 => "110101100111",
    3432 => "110101101000",
    3433 => "110101101001",
    3434 => "110101101010",
    3435 => "110101101011",
    3436 => "110101101100",
    3437 => "110101101101",
    3438 => "110101101110",
    3439 => "110101101111",
    3440 => "110101110000",
    3441 => "110101110001",
    3442 => "110101110010",
    3443 => "110101110011",
    3444 => "110101110100",
    3445 => "110101110101",
    3446 => "110101110110",
    3447 => "110101110111",
    3448 => "110101111000",
    3449 => "110101111001",
    3450 => "110101111010",
    3451 => "110101111011",
    3452 => "110101111100",
    3453 => "110101111101",
    3454 => "110101111110",
    3455 => "110101111111",
    3456 => "110110000000",
    3457 => "110110000001",
    3458 => "110110000010",
    3459 => "110110000011",
    3460 => "110110000100",
    3461 => "110110000101",
    3462 => "110110000110",
    3463 => "110110000111",
    3464 => "110110001000",
    3465 => "110110001001",
    3466 => "110110001010",
    3467 => "110110001011",
    3468 => "110110001100",
    3469 => "110110001101",
    3470 => "110110001110",
    3471 => "110110001111",
    3472 => "110110010000",
    3473 => "110110010001",
    3474 => "110110010010",
    3475 => "110110010011",
    3476 => "110110010100",
    3477 => "110110010101",
    3478 => "110110010110",
    3479 => "110110010111",
    3480 => "110110011000",
    3481 => "110110011001",
    3482 => "110110011010",
    3483 => "110110011011",
    3484 => "110110011100",
    3485 => "110110011101",
    3486 => "110110011110",
    3487 => "110110011111",
    3488 => "110110100000",
    3489 => "110110100001",
    3490 => "110110100010",
    3491 => "110110100011",
    3492 => "110110100100",
    3493 => "110110100101",
    3494 => "110110100110",
    3495 => "110110100111",
    3496 => "110110101000",
    3497 => "110110101001",
    3498 => "110110101010",
    3499 => "110110101011",
    3500 => "110110101100",
    3501 => "110110101101",
    3502 => "110110101110",
    3503 => "110110101111",
    3504 => "110110110000",
    3505 => "110110110001",
    3506 => "110110110010",
    3507 => "110110110011",
    3508 => "110110110100",
    3509 => "110110110101",
    3510 => "110110110110",
    3511 => "110110110111",
    3512 => "110110111000",
    3513 => "110110111001",
    3514 => "110110111010",
    3515 => "110110111011",
    3516 => "110110111100",
    3517 => "110110111101",
    3518 => "110110111110",
    3519 => "110110111111",
    3520 => "110111000000",
    3521 => "110111000001",
    3522 => "110111000010",
    3523 => "110111000011",
    3524 => "110111000100",
    3525 => "110111000101",
    3526 => "110111000110",
    3527 => "110111000111",
    3528 => "110111001000",
    3529 => "110111001001",
    3530 => "110111001010",
    3531 => "110111001011",
    3532 => "110111001100",
    3533 => "110111001101",
    3534 => "110111001110",
    3535 => "110111001111",
    3536 => "110111010000",
    3537 => "110111010001",
    3538 => "110111010010",
    3539 => "110111010011",
    3540 => "110111010100",
    3541 => "110111010101",
    3542 => "110111010110",
    3543 => "110111010111",
    3544 => "110111011000",
    3545 => "110111011001",
    3546 => "110111011010",
    3547 => "110111011011",
    3548 => "110111011100",
    3549 => "110111011101",
    3550 => "110111011110",
    3551 => "110111011111",
    3552 => "110111100000",
    3553 => "110111100001",
    3554 => "110111100010",
    3555 => "110111100011",
    3556 => "110111100100",
    3557 => "110111100101",
    3558 => "110111100110",
    3559 => "110111100111",
    3560 => "110111101000",
    3561 => "110111101001",
    3562 => "110111101010",
    3563 => "110111101011",
    3564 => "110111101100",
    3565 => "110111101101",
    3566 => "110111101110",
    3567 => "110111101111",
    3568 => "110111110000",
    3569 => "110111110001",
    3570 => "110111110010",
    3571 => "110111110011",
    3572 => "110111110100",
    3573 => "110111110101",
    3574 => "110111110110",
    3575 => "110111110111",
    3576 => "110111111000",
    3577 => "110111111001",
    3578 => "110111111010",
    3579 => "110111111011",
    3580 => "110111111100",
    3581 => "110111111101",
    3582 => "110111111110",
    3583 => "110111111111",
    3584 => "111000000000",
    3585 => "111000000001",
    3586 => "111000000010",
    3587 => "111000000011",
    3588 => "111000000100",
    3589 => "111000000101",
    3590 => "111000000110",
    3591 => "111000000111",
    3592 => "111000001000",
    3593 => "111000001001",
    3594 => "111000001010",
    3595 => "111000001011",
    3596 => "111000001100",
    3597 => "111000001101",
    3598 => "111000001110",
    3599 => "111000001111",
    3600 => "111000010000",
    3601 => "111000010001",
    3602 => "111000010010",
    3603 => "111000010011",
    3604 => "111000010100",
    3605 => "111000010101",
    3606 => "111000010110",
    3607 => "111000010111",
    3608 => "111000011000",
    3609 => "111000011001",
    3610 => "111000011010",
    3611 => "111000011011",
    3612 => "111000011100",
    3613 => "111000011101",
    3614 => "111000011110",
    3615 => "111000011111",
    3616 => "111000100000",
    3617 => "111000100001",
    3618 => "111000100010",
    3619 => "111000100011",
    3620 => "111000100100",
    3621 => "111000100101",
    3622 => "111000100110",
    3623 => "111000100111",
    3624 => "111000101000",
    3625 => "111000101001",
    3626 => "111000101010",
    3627 => "111000101011",
    3628 => "111000101100",
    3629 => "111000101101",
    3630 => "111000101110",
    3631 => "111000101111",
    3632 => "111000110000",
    3633 => "111000110001",
    3634 => "111000110010",
    3635 => "111000110011",
    3636 => "111000110100",
    3637 => "111000110101",
    3638 => "111000110110",
    3639 => "111000110111",
    3640 => "111000111000",
    3641 => "111000111001",
    3642 => "111000111010",
    3643 => "111000111011",
    3644 => "111000111100",
    3645 => "111000111101",
    3646 => "111000111110",
    3647 => "111000111111",
    3648 => "111001000000",
    3649 => "111001000001",
    3650 => "111001000010",
    3651 => "111001000011",
    3652 => "111001000100",
    3653 => "111001000101",
    3654 => "111001000110",
    3655 => "111001000111",
    3656 => "111001001000",
    3657 => "111001001001",
    3658 => "111001001010",
    3659 => "111001001011",
    3660 => "111001001100",
    3661 => "111001001101",
    3662 => "111001001110",
    3663 => "111001001111",
    3664 => "111001010000",
    3665 => "111001010001",
    3666 => "111001010010",
    3667 => "111001010011",
    3668 => "111001010100",
    3669 => "111001010101",
    3670 => "111001010110",
    3671 => "111001010111",
    3672 => "111001011000",
    3673 => "111001011001",
    3674 => "111001011010",
    3675 => "111001011011",
    3676 => "111001011100",
    3677 => "111001011101",
    3678 => "111001011110",
    3679 => "111001011111",
    3680 => "111001100000",
    3681 => "111001100001",
    3682 => "111001100010",
    3683 => "111001100011",
    3684 => "111001100100",
    3685 => "111001100101",
    3686 => "111001100110",
    3687 => "111001100111",
    3688 => "111001101000",
    3689 => "111001101001",
    3690 => "111001101010",
    3691 => "111001101011",
    3692 => "111001101100",
    3693 => "111001101101",
    3694 => "111001101110",
    3695 => "111001101111",
    3696 => "111001110000",
    3697 => "111001110001",
    3698 => "111001110010",
    3699 => "111001110011",
    3700 => "111001110100",
    3701 => "111001110101",
    3702 => "111001110110",
    3703 => "111001110111",
    3704 => "111001111000",
    3705 => "111001111001",
    3706 => "111001111010",
    3707 => "111001111011",
    3708 => "111001111100",
    3709 => "111001111101",
    3710 => "111001111110",
    3711 => "111001111111",
    3712 => "111010000000",
    3713 => "111010000001",
    3714 => "111010000010",
    3715 => "111010000011",
    3716 => "111010000100",
    3717 => "111010000101",
    3718 => "111010000110",
    3719 => "111010000111",
    3720 => "111010001000",
    3721 => "111010001001",
    3722 => "111010001010",
    3723 => "111010001011",
    3724 => "111010001100",
    3725 => "111010001101",
    3726 => "111010001110",
    3727 => "111010001111",
    3728 => "111010010000",
    3729 => "111010010001",
    3730 => "111010010010",
    3731 => "111010010011",
    3732 => "111010010100",
    3733 => "111010010101",
    3734 => "111010010110",
    3735 => "111010010111",
    3736 => "111010011000",
    3737 => "111010011001",
    3738 => "111010011010",
    3739 => "111010011011",
    3740 => "111010011100",
    3741 => "111010011101",
    3742 => "111010011110",
    3743 => "111010011111",
    3744 => "111010100000",
    3745 => "111010100001",
    3746 => "111010100010",
    3747 => "111010100011",
    3748 => "111010100100",
    3749 => "111010100101",
    3750 => "111010100110",
    3751 => "111010100111",
    3752 => "111010101000",
    3753 => "111010101001",
    3754 => "111010101010",
    3755 => "111010101011",
    3756 => "111010101100",
    3757 => "111010101101",
    3758 => "111010101110",
    3759 => "111010101111",
    3760 => "111010110000",
    3761 => "111010110001",
    3762 => "111010110010",
    3763 => "111010110011",
    3764 => "111010110100",
    3765 => "111010110101",
    3766 => "111010110110",
    3767 => "111010110111",
    3768 => "111010111000",
    3769 => "111010111001",
    3770 => "111010111010",
    3771 => "111010111011",
    3772 => "111010111100",
    3773 => "111010111101",
    3774 => "111010111110",
    3775 => "111010111111",
    3776 => "111011000000",
    3777 => "111011000001",
    3778 => "111011000010",
    3779 => "111011000011",
    3780 => "111011000100",
    3781 => "111011000101",
    3782 => "111011000110",
    3783 => "111011000111",
    3784 => "111011001000",
    3785 => "111011001001",
    3786 => "111011001010",
    3787 => "111011001011",
    3788 => "111011001100",
    3789 => "111011001101",
    3790 => "111011001110",
    3791 => "111011001111",
    3792 => "111011010000",
    3793 => "111011010001",
    3794 => "111011010010",
    3795 => "111011010011",
    3796 => "111011010100",
    3797 => "111011010101",
    3798 => "111011010110",
    3799 => "111011010111",
    3800 => "111011011000",
    3801 => "111011011001",
    3802 => "111011011010",
    3803 => "111011011011",
    3804 => "111011011100",
    3805 => "111011011101",
    3806 => "111011011110",
    3807 => "111011011111",
    3808 => "111011100000",
    3809 => "111011100001",
    3810 => "111011100010",
    3811 => "111011100011",
    3812 => "111011100100",
    3813 => "111011100101",
    3814 => "111011100110",
    3815 => "111011100111",
    3816 => "111011101000",
    3817 => "111011101001",
    3818 => "111011101010",
    3819 => "111011101011",
    3820 => "111011101100",
    3821 => "111011101101",
    3822 => "111011101110",
    3823 => "111011101111",
    3824 => "111011110000",
    3825 => "111011110001",
    3826 => "111011110010",
    3827 => "111011110011",
    3828 => "111011110100",
    3829 => "111011110101",
    3830 => "111011110110",
    3831 => "111011110111",
    3832 => "111011111000",
    3833 => "111011111001",
    3834 => "111011111010",
    3835 => "111011111011",
    3836 => "111011111100",
    3837 => "111011111101",
    3838 => "111011111110",
    3839 => "111011111111",
    3840 => "111100000000",
    3841 => "111100000001",
    3842 => "111100000010",
    3843 => "111100000011",
    3844 => "111100000100",
    3845 => "111100000101",
    3846 => "111100000110",
    3847 => "111100000111",
    3848 => "111100001000",
    3849 => "111100001001",
    3850 => "111100001010",
    3851 => "111100001011",
    3852 => "111100001100",
    3853 => "111100001101",
    3854 => "111100001110",
    3855 => "111100001111",
    3856 => "111100010000",
    3857 => "111100010001",
    3858 => "111100010010",
    3859 => "111100010011",
    3860 => "111100010100",
    3861 => "111100010101",
    3862 => "111100010110",
    3863 => "111100010111",
    3864 => "111100011000",
    3865 => "111100011001",
    3866 => "111100011010",
    3867 => "111100011011",
    3868 => "111100011100",
    3869 => "111100011101",
    3870 => "111100011110",
    3871 => "111100011111",
    3872 => "111100100000",
    3873 => "111100100001",
    3874 => "111100100010",
    3875 => "111100100011",
    3876 => "111100100100",
    3877 => "111100100101",
    3878 => "111100100110",
    3879 => "111100100111",
    3880 => "111100101000",
    3881 => "111100101001",
    3882 => "111100101010",
    3883 => "111100101011",
    3884 => "111100101100",
    3885 => "111100101101",
    3886 => "111100101110",
    3887 => "111100101111",
    3888 => "111100110000",
    3889 => "111100110001",
    3890 => "111100110010",
    3891 => "111100110011",
    3892 => "111100110100",
    3893 => "111100110101",
    3894 => "111100110110",
    3895 => "111100110111",
    3896 => "111100111000",
    3897 => "111100111001",
    3898 => "111100111010",
    3899 => "111100111011",
    3900 => "111100111100",
    3901 => "111100111101",
    3902 => "111100111110",
    3903 => "111100111111",
    3904 => "111101000000",
    3905 => "111101000001",
    3906 => "111101000010",
    3907 => "111101000011",
    3908 => "111101000100",
    3909 => "111101000101",
    3910 => "111101000110",
    3911 => "111101000111",
    3912 => "111101001000",
    3913 => "111101001001",
    3914 => "111101001010",
    3915 => "111101001011",
    3916 => "111101001100",
    3917 => "111101001101",
    3918 => "111101001110",
    3919 => "111101001111",
    3920 => "111101010000",
    3921 => "111101010001",
    3922 => "111101010010",
    3923 => "111101010011",
    3924 => "111101010100",
    3925 => "111101010101",
    3926 => "111101010110",
    3927 => "111101010111",
    3928 => "111101011000",
    3929 => "111101011001",
    3930 => "111101011010",
    3931 => "111101011011",
    3932 => "111101011100",
    3933 => "111101011101",
    3934 => "111101011110",
    3935 => "111101011111",
    3936 => "111101100000",
    3937 => "111101100001",
    3938 => "111101100010",
    3939 => "111101100011",
    3940 => "111101100100",
    3941 => "111101100101",
    3942 => "111101100110",
    3943 => "111101100111",
    3944 => "111101101000",
    3945 => "111101101001",
    3946 => "111101101010",
    3947 => "111101101011",
    3948 => "111101101100",
    3949 => "111101101101",
    3950 => "111101101110",
    3951 => "111101101111",
    3952 => "111101110000",
    3953 => "111101110001",
    3954 => "111101110010",
    3955 => "111101110011",
    3956 => "111101110100",
    3957 => "111101110101",
    3958 => "111101110110",
    3959 => "111101110111",
    3960 => "111101111000",
    3961 => "111101111001",
    3962 => "111101111010",
    3963 => "111101111011",
    3964 => "111101111100",
    3965 => "111101111101",
    3966 => "111101111110",
    3967 => "111101111111",
    3968 => "111110000000",
    3969 => "111110000001",
    3970 => "111110000010",
    3971 => "111110000011",
    3972 => "111110000100",
    3973 => "111110000101",
    3974 => "111110000110",
    3975 => "111110000111",
    3976 => "111110001000",
    3977 => "111110001001",
    3978 => "111110001010",
    3979 => "111110001011",
    3980 => "111110001100",
    3981 => "111110001101",
    3982 => "111110001110",
    3983 => "111110001111",
    3984 => "111110010000",
    3985 => "111110010001",
    3986 => "111110010010",
    3987 => "111110010011",
    3988 => "111110010100",
    3989 => "111110010101",
    3990 => "111110010110",
    3991 => "111110010111",
    3992 => "111110011000",
    3993 => "111110011001",
    3994 => "111110011010",
    3995 => "111110011011",
    3996 => "111110011100",
    3997 => "111110011101",
    3998 => "111110011110",
    3999 => "111110011111",
    4000 => "111110100000",
    4001 => "111110100001",
    4002 => "111110100010",
    4003 => "111110100011",
    4004 => "111110100100",
    4005 => "111110100101",
    4006 => "111110100110",
    4007 => "111110100111",
    4008 => "111110101000",
    4009 => "111110101001",
    4010 => "111110101010",
    4011 => "111110101011",
    4012 => "111110101100",
    4013 => "111110101101",
    4014 => "111110101110",
    4015 => "111110101111",
    4016 => "111110110000",
    4017 => "111110110001",
    4018 => "111110110010",
    4019 => "111110110011",
    4020 => "111110110100",
    4021 => "111110110101",
    4022 => "111110110110",
    4023 => "111110110111",
    4024 => "111110111000",
    4025 => "111110111001",
    4026 => "111110111010",
    4027 => "111110111011",
    4028 => "111110111100",
    4029 => "111110111101",
    4030 => "111110111110",
    4031 => "111110111111",
    4032 => "111111000000",
    4033 => "111111000001",
    4034 => "111111000010",
    4035 => "111111000011",
    4036 => "111111000100",
    4037 => "111111000101",
    4038 => "111111000110",
    4039 => "111111000111",
    4040 => "111111001000",
    4041 => "111111001001",
    4042 => "111111001010",
    4043 => "111111001011",
    4044 => "111111001100",
    4045 => "111111001101",
    4046 => "111111001110",
    4047 => "111111001111",
    4048 => "111111010000",
    4049 => "111111010001",
    4050 => "111111010010",
    4051 => "111111010011",
    4052 => "111111010100",
    4053 => "111111010101",
    4054 => "111111010110",
    4055 => "111111010111",
    4056 => "111111011000",
    4057 => "111111011001",
    4058 => "111111011010",
    4059 => "111111011011",
    4060 => "111111011100",
    4061 => "111111011101",
    4062 => "111111011110",
    4063 => "111111011111",
    4064 => "111111100000",
    4065 => "111111100001",
    4066 => "111111100010",
    4067 => "111111100011",
    4068 => "111111100100",
    4069 => "111111100101",
    4070 => "111111100110",
    4071 => "111111100111",
    4072 => "111111101000",
    4073 => "111111101001",
    4074 => "111111101010",
    4075 => "111111101011",
    4076 => "111111101100",
    4077 => "111111101101",
    4078 => "111111101110",
    4079 => "111111101111",
    4080 => "111111110000",
    4081 => "111111110001",
    4082 => "111111110010",
    4083 => "111111110011",
    4084 => "111111110100",
    4085 => "111111110101",
    4086 => "111111110110",
    4087 => "111111110111",
    4088 => "111111111000",
    4089 => "111111111001",
    4090 => "111111111010",
    4091 => "111111111011",
    4092 => "111111111100",
    4093 => "111111111101",
    4094 => "111111111110",
    4095 => "111111111110");
begin
 process (address)
 begin
  case address is
     when "000000000000" => data <= saw_rom(0);
     when "000000000001" => data <= saw_rom(1);
     when "000000000010" => data <= saw_rom(2);
     when "000000000011" => data <= saw_rom(3);
     when "000000000100" => data <= saw_rom(4);
     when "000000000101" => data <= saw_rom(5);
     when "000000000110" => data <= saw_rom(6);
     when "000000000111" => data <= saw_rom(7);
     when "000000001000" => data <= saw_rom(8);
     when "000000001001" => data <= saw_rom(9);
     when "000000001010" => data <= saw_rom(10);
     when "000000001011" => data <= saw_rom(11);
     when "000000001100" => data <= saw_rom(12);
     when "000000001101" => data <= saw_rom(13);
     when "000000001110" => data <= saw_rom(14);
     when "000000001111" => data <= saw_rom(15);
     when "000000010000" => data <= saw_rom(16);
     when "000000010001" => data <= saw_rom(17);
     when "000000010010" => data <= saw_rom(18);
     when "000000010011" => data <= saw_rom(19);
     when "000000010100" => data <= saw_rom(20);
     when "000000010101" => data <= saw_rom(21);
     when "000000010110" => data <= saw_rom(22);
     when "000000010111" => data <= saw_rom(23);
     when "000000011000" => data <= saw_rom(24);
     when "000000011001" => data <= saw_rom(25);
     when "000000011010" => data <= saw_rom(26);
     when "000000011011" => data <= saw_rom(27);
     when "000000011100" => data <= saw_rom(28);
     when "000000011101" => data <= saw_rom(29);
     when "000000011110" => data <= saw_rom(30);
     when "000000011111" => data <= saw_rom(31);
     when "000000100000" => data <= saw_rom(32);
     when "000000100001" => data <= saw_rom(33);
     when "000000100010" => data <= saw_rom(34);
     when "000000100011" => data <= saw_rom(35);
     when "000000100100" => data <= saw_rom(36);
     when "000000100101" => data <= saw_rom(37);
     when "000000100110" => data <= saw_rom(38);
     when "000000100111" => data <= saw_rom(39);
     when "000000101000" => data <= saw_rom(40);
     when "000000101001" => data <= saw_rom(41);
     when "000000101010" => data <= saw_rom(42);
     when "000000101011" => data <= saw_rom(43);
     when "000000101100" => data <= saw_rom(44);
     when "000000101101" => data <= saw_rom(45);
     when "000000101110" => data <= saw_rom(46);
     when "000000101111" => data <= saw_rom(47);
     when "000000110000" => data <= saw_rom(48);
     when "000000110001" => data <= saw_rom(49);
     when "000000110010" => data <= saw_rom(50);
     when "000000110011" => data <= saw_rom(51);
     when "000000110100" => data <= saw_rom(52);
     when "000000110101" => data <= saw_rom(53);
     when "000000110110" => data <= saw_rom(54);
     when "000000110111" => data <= saw_rom(55);
     when "000000111000" => data <= saw_rom(56);
     when "000000111001" => data <= saw_rom(57);
     when "000000111010" => data <= saw_rom(58);
     when "000000111011" => data <= saw_rom(59);
     when "000000111100" => data <= saw_rom(60);
     when "000000111101" => data <= saw_rom(61);
     when "000000111110" => data <= saw_rom(62);
     when "000000111111" => data <= saw_rom(63);
     when "000001000000" => data <= saw_rom(64);
     when "000001000001" => data <= saw_rom(65);
     when "000001000010" => data <= saw_rom(66);
     when "000001000011" => data <= saw_rom(67);
     when "000001000100" => data <= saw_rom(68);
     when "000001000101" => data <= saw_rom(69);
     when "000001000110" => data <= saw_rom(70);
     when "000001000111" => data <= saw_rom(71);
     when "000001001000" => data <= saw_rom(72);
     when "000001001001" => data <= saw_rom(73);
     when "000001001010" => data <= saw_rom(74);
     when "000001001011" => data <= saw_rom(75);
     when "000001001100" => data <= saw_rom(76);
     when "000001001101" => data <= saw_rom(77);
     when "000001001110" => data <= saw_rom(78);
     when "000001001111" => data <= saw_rom(79);
     when "000001010000" => data <= saw_rom(80);
     when "000001010001" => data <= saw_rom(81);
     when "000001010010" => data <= saw_rom(82);
     when "000001010011" => data <= saw_rom(83);
     when "000001010100" => data <= saw_rom(84);
     when "000001010101" => data <= saw_rom(85);
     when "000001010110" => data <= saw_rom(86);
     when "000001010111" => data <= saw_rom(87);
     when "000001011000" => data <= saw_rom(88);
     when "000001011001" => data <= saw_rom(89);
     when "000001011010" => data <= saw_rom(90);
     when "000001011011" => data <= saw_rom(91);
     when "000001011100" => data <= saw_rom(92);
     when "000001011101" => data <= saw_rom(93);
     when "000001011110" => data <= saw_rom(94);
     when "000001011111" => data <= saw_rom(95);
     when "000001100000" => data <= saw_rom(96);
     when "000001100001" => data <= saw_rom(97);
     when "000001100010" => data <= saw_rom(98);
     when "000001100011" => data <= saw_rom(99);
     when "000001100100" => data <= saw_rom(100);
     when "000001100101" => data <= saw_rom(101);
     when "000001100110" => data <= saw_rom(102);
     when "000001100111" => data <= saw_rom(103);
     when "000001101000" => data <= saw_rom(104);
     when "000001101001" => data <= saw_rom(105);
     when "000001101010" => data <= saw_rom(106);
     when "000001101011" => data <= saw_rom(107);
     when "000001101100" => data <= saw_rom(108);
     when "000001101101" => data <= saw_rom(109);
     when "000001101110" => data <= saw_rom(110);
     when "000001101111" => data <= saw_rom(111);
     when "000001110000" => data <= saw_rom(112);
     when "000001110001" => data <= saw_rom(113);
     when "000001110010" => data <= saw_rom(114);
     when "000001110011" => data <= saw_rom(115);
     when "000001110100" => data <= saw_rom(116);
     when "000001110101" => data <= saw_rom(117);
     when "000001110110" => data <= saw_rom(118);
     when "000001110111" => data <= saw_rom(119);
     when "000001111000" => data <= saw_rom(120);
     when "000001111001" => data <= saw_rom(121);
     when "000001111010" => data <= saw_rom(122);
     when "000001111011" => data <= saw_rom(123);
     when "000001111100" => data <= saw_rom(124);
     when "000001111101" => data <= saw_rom(125);
     when "000001111110" => data <= saw_rom(126);
     when "000001111111" => data <= saw_rom(127);
     when "000010000000" => data <= saw_rom(128);
     when "000010000001" => data <= saw_rom(129);
     when "000010000010" => data <= saw_rom(130);
     when "000010000011" => data <= saw_rom(131);
     when "000010000100" => data <= saw_rom(132);
     when "000010000101" => data <= saw_rom(133);
     when "000010000110" => data <= saw_rom(134);
     when "000010000111" => data <= saw_rom(135);
     when "000010001000" => data <= saw_rom(136);
     when "000010001001" => data <= saw_rom(137);
     when "000010001010" => data <= saw_rom(138);
     when "000010001011" => data <= saw_rom(139);
     when "000010001100" => data <= saw_rom(140);
     when "000010001101" => data <= saw_rom(141);
     when "000010001110" => data <= saw_rom(142);
     when "000010001111" => data <= saw_rom(143);
     when "000010010000" => data <= saw_rom(144);
     when "000010010001" => data <= saw_rom(145);
     when "000010010010" => data <= saw_rom(146);
     when "000010010011" => data <= saw_rom(147);
     when "000010010100" => data <= saw_rom(148);
     when "000010010101" => data <= saw_rom(149);
     when "000010010110" => data <= saw_rom(150);
     when "000010010111" => data <= saw_rom(151);
     when "000010011000" => data <= saw_rom(152);
     when "000010011001" => data <= saw_rom(153);
     when "000010011010" => data <= saw_rom(154);
     when "000010011011" => data <= saw_rom(155);
     when "000010011100" => data <= saw_rom(156);
     when "000010011101" => data <= saw_rom(157);
     when "000010011110" => data <= saw_rom(158);
     when "000010011111" => data <= saw_rom(159);
     when "000010100000" => data <= saw_rom(160);
     when "000010100001" => data <= saw_rom(161);
     when "000010100010" => data <= saw_rom(162);
     when "000010100011" => data <= saw_rom(163);
     when "000010100100" => data <= saw_rom(164);
     when "000010100101" => data <= saw_rom(165);
     when "000010100110" => data <= saw_rom(166);
     when "000010100111" => data <= saw_rom(167);
     when "000010101000" => data <= saw_rom(168);
     when "000010101001" => data <= saw_rom(169);
     when "000010101010" => data <= saw_rom(170);
     when "000010101011" => data <= saw_rom(171);
     when "000010101100" => data <= saw_rom(172);
     when "000010101101" => data <= saw_rom(173);
     when "000010101110" => data <= saw_rom(174);
     when "000010101111" => data <= saw_rom(175);
     when "000010110000" => data <= saw_rom(176);
     when "000010110001" => data <= saw_rom(177);
     when "000010110010" => data <= saw_rom(178);
     when "000010110011" => data <= saw_rom(179);
     when "000010110100" => data <= saw_rom(180);
     when "000010110101" => data <= saw_rom(181);
     when "000010110110" => data <= saw_rom(182);
     when "000010110111" => data <= saw_rom(183);
     when "000010111000" => data <= saw_rom(184);
     when "000010111001" => data <= saw_rom(185);
     when "000010111010" => data <= saw_rom(186);
     when "000010111011" => data <= saw_rom(187);
     when "000010111100" => data <= saw_rom(188);
     when "000010111101" => data <= saw_rom(189);
     when "000010111110" => data <= saw_rom(190);
     when "000010111111" => data <= saw_rom(191);
     when "000011000000" => data <= saw_rom(192);
     when "000011000001" => data <= saw_rom(193);
     when "000011000010" => data <= saw_rom(194);
     when "000011000011" => data <= saw_rom(195);
     when "000011000100" => data <= saw_rom(196);
     when "000011000101" => data <= saw_rom(197);
     when "000011000110" => data <= saw_rom(198);
     when "000011000111" => data <= saw_rom(199);
     when "000011001000" => data <= saw_rom(200);
     when "000011001001" => data <= saw_rom(201);
     when "000011001010" => data <= saw_rom(202);
     when "000011001011" => data <= saw_rom(203);
     when "000011001100" => data <= saw_rom(204);
     when "000011001101" => data <= saw_rom(205);
     when "000011001110" => data <= saw_rom(206);
     when "000011001111" => data <= saw_rom(207);
     when "000011010000" => data <= saw_rom(208);
     when "000011010001" => data <= saw_rom(209);
     when "000011010010" => data <= saw_rom(210);
     when "000011010011" => data <= saw_rom(211);
     when "000011010100" => data <= saw_rom(212);
     when "000011010101" => data <= saw_rom(213);
     when "000011010110" => data <= saw_rom(214);
     when "000011010111" => data <= saw_rom(215);
     when "000011011000" => data <= saw_rom(216);
     when "000011011001" => data <= saw_rom(217);
     when "000011011010" => data <= saw_rom(218);
     when "000011011011" => data <= saw_rom(219);
     when "000011011100" => data <= saw_rom(220);
     when "000011011101" => data <= saw_rom(221);
     when "000011011110" => data <= saw_rom(222);
     when "000011011111" => data <= saw_rom(223);
     when "000011100000" => data <= saw_rom(224);
     when "000011100001" => data <= saw_rom(225);
     when "000011100010" => data <= saw_rom(226);
     when "000011100011" => data <= saw_rom(227);
     when "000011100100" => data <= saw_rom(228);
     when "000011100101" => data <= saw_rom(229);
     when "000011100110" => data <= saw_rom(230);
     when "000011100111" => data <= saw_rom(231);
     when "000011101000" => data <= saw_rom(232);
     when "000011101001" => data <= saw_rom(233);
     when "000011101010" => data <= saw_rom(234);
     when "000011101011" => data <= saw_rom(235);
     when "000011101100" => data <= saw_rom(236);
     when "000011101101" => data <= saw_rom(237);
     when "000011101110" => data <= saw_rom(238);
     when "000011101111" => data <= saw_rom(239);
     when "000011110000" => data <= saw_rom(240);
     when "000011110001" => data <= saw_rom(241);
     when "000011110010" => data <= saw_rom(242);
     when "000011110011" => data <= saw_rom(243);
     when "000011110100" => data <= saw_rom(244);
     when "000011110101" => data <= saw_rom(245);
     when "000011110110" => data <= saw_rom(246);
     when "000011110111" => data <= saw_rom(247);
     when "000011111000" => data <= saw_rom(248);
     when "000011111001" => data <= saw_rom(249);
     when "000011111010" => data <= saw_rom(250);
     when "000011111011" => data <= saw_rom(251);
     when "000011111100" => data <= saw_rom(252);
     when "000011111101" => data <= saw_rom(253);
     when "000011111110" => data <= saw_rom(254);
     when "000011111111" => data <= saw_rom(255);
     when "000100000000" => data <= saw_rom(256);
     when "000100000001" => data <= saw_rom(257);
     when "000100000010" => data <= saw_rom(258);
     when "000100000011" => data <= saw_rom(259);
     when "000100000100" => data <= saw_rom(260);
     when "000100000101" => data <= saw_rom(261);
     when "000100000110" => data <= saw_rom(262);
     when "000100000111" => data <= saw_rom(263);
     when "000100001000" => data <= saw_rom(264);
     when "000100001001" => data <= saw_rom(265);
     when "000100001010" => data <= saw_rom(266);
     when "000100001011" => data <= saw_rom(267);
     when "000100001100" => data <= saw_rom(268);
     when "000100001101" => data <= saw_rom(269);
     when "000100001110" => data <= saw_rom(270);
     when "000100001111" => data <= saw_rom(271);
     when "000100010000" => data <= saw_rom(272);
     when "000100010001" => data <= saw_rom(273);
     when "000100010010" => data <= saw_rom(274);
     when "000100010011" => data <= saw_rom(275);
     when "000100010100" => data <= saw_rom(276);
     when "000100010101" => data <= saw_rom(277);
     when "000100010110" => data <= saw_rom(278);
     when "000100010111" => data <= saw_rom(279);
     when "000100011000" => data <= saw_rom(280);
     when "000100011001" => data <= saw_rom(281);
     when "000100011010" => data <= saw_rom(282);
     when "000100011011" => data <= saw_rom(283);
     when "000100011100" => data <= saw_rom(284);
     when "000100011101" => data <= saw_rom(285);
     when "000100011110" => data <= saw_rom(286);
     when "000100011111" => data <= saw_rom(287);
     when "000100100000" => data <= saw_rom(288);
     when "000100100001" => data <= saw_rom(289);
     when "000100100010" => data <= saw_rom(290);
     when "000100100011" => data <= saw_rom(291);
     when "000100100100" => data <= saw_rom(292);
     when "000100100101" => data <= saw_rom(293);
     when "000100100110" => data <= saw_rom(294);
     when "000100100111" => data <= saw_rom(295);
     when "000100101000" => data <= saw_rom(296);
     when "000100101001" => data <= saw_rom(297);
     when "000100101010" => data <= saw_rom(298);
     when "000100101011" => data <= saw_rom(299);
     when "000100101100" => data <= saw_rom(300);
     when "000100101101" => data <= saw_rom(301);
     when "000100101110" => data <= saw_rom(302);
     when "000100101111" => data <= saw_rom(303);
     when "000100110000" => data <= saw_rom(304);
     when "000100110001" => data <= saw_rom(305);
     when "000100110010" => data <= saw_rom(306);
     when "000100110011" => data <= saw_rom(307);
     when "000100110100" => data <= saw_rom(308);
     when "000100110101" => data <= saw_rom(309);
     when "000100110110" => data <= saw_rom(310);
     when "000100110111" => data <= saw_rom(311);
     when "000100111000" => data <= saw_rom(312);
     when "000100111001" => data <= saw_rom(313);
     when "000100111010" => data <= saw_rom(314);
     when "000100111011" => data <= saw_rom(315);
     when "000100111100" => data <= saw_rom(316);
     when "000100111101" => data <= saw_rom(317);
     when "000100111110" => data <= saw_rom(318);
     when "000100111111" => data <= saw_rom(319);
     when "000101000000" => data <= saw_rom(320);
     when "000101000001" => data <= saw_rom(321);
     when "000101000010" => data <= saw_rom(322);
     when "000101000011" => data <= saw_rom(323);
     when "000101000100" => data <= saw_rom(324);
     when "000101000101" => data <= saw_rom(325);
     when "000101000110" => data <= saw_rom(326);
     when "000101000111" => data <= saw_rom(327);
     when "000101001000" => data <= saw_rom(328);
     when "000101001001" => data <= saw_rom(329);
     when "000101001010" => data <= saw_rom(330);
     when "000101001011" => data <= saw_rom(331);
     when "000101001100" => data <= saw_rom(332);
     when "000101001101" => data <= saw_rom(333);
     when "000101001110" => data <= saw_rom(334);
     when "000101001111" => data <= saw_rom(335);
     when "000101010000" => data <= saw_rom(336);
     when "000101010001" => data <= saw_rom(337);
     when "000101010010" => data <= saw_rom(338);
     when "000101010011" => data <= saw_rom(339);
     when "000101010100" => data <= saw_rom(340);
     when "000101010101" => data <= saw_rom(341);
     when "000101010110" => data <= saw_rom(342);
     when "000101010111" => data <= saw_rom(343);
     when "000101011000" => data <= saw_rom(344);
     when "000101011001" => data <= saw_rom(345);
     when "000101011010" => data <= saw_rom(346);
     when "000101011011" => data <= saw_rom(347);
     when "000101011100" => data <= saw_rom(348);
     when "000101011101" => data <= saw_rom(349);
     when "000101011110" => data <= saw_rom(350);
     when "000101011111" => data <= saw_rom(351);
     when "000101100000" => data <= saw_rom(352);
     when "000101100001" => data <= saw_rom(353);
     when "000101100010" => data <= saw_rom(354);
     when "000101100011" => data <= saw_rom(355);
     when "000101100100" => data <= saw_rom(356);
     when "000101100101" => data <= saw_rom(357);
     when "000101100110" => data <= saw_rom(358);
     when "000101100111" => data <= saw_rom(359);
     when "000101101000" => data <= saw_rom(360);
     when "000101101001" => data <= saw_rom(361);
     when "000101101010" => data <= saw_rom(362);
     when "000101101011" => data <= saw_rom(363);
     when "000101101100" => data <= saw_rom(364);
     when "000101101101" => data <= saw_rom(365);
     when "000101101110" => data <= saw_rom(366);
     when "000101101111" => data <= saw_rom(367);
     when "000101110000" => data <= saw_rom(368);
     when "000101110001" => data <= saw_rom(369);
     when "000101110010" => data <= saw_rom(370);
     when "000101110011" => data <= saw_rom(371);
     when "000101110100" => data <= saw_rom(372);
     when "000101110101" => data <= saw_rom(373);
     when "000101110110" => data <= saw_rom(374);
     when "000101110111" => data <= saw_rom(375);
     when "000101111000" => data <= saw_rom(376);
     when "000101111001" => data <= saw_rom(377);
     when "000101111010" => data <= saw_rom(378);
     when "000101111011" => data <= saw_rom(379);
     when "000101111100" => data <= saw_rom(380);
     when "000101111101" => data <= saw_rom(381);
     when "000101111110" => data <= saw_rom(382);
     when "000101111111" => data <= saw_rom(383);
     when "000110000000" => data <= saw_rom(384);
     when "000110000001" => data <= saw_rom(385);
     when "000110000010" => data <= saw_rom(386);
     when "000110000011" => data <= saw_rom(387);
     when "000110000100" => data <= saw_rom(388);
     when "000110000101" => data <= saw_rom(389);
     when "000110000110" => data <= saw_rom(390);
     when "000110000111" => data <= saw_rom(391);
     when "000110001000" => data <= saw_rom(392);
     when "000110001001" => data <= saw_rom(393);
     when "000110001010" => data <= saw_rom(394);
     when "000110001011" => data <= saw_rom(395);
     when "000110001100" => data <= saw_rom(396);
     when "000110001101" => data <= saw_rom(397);
     when "000110001110" => data <= saw_rom(398);
     when "000110001111" => data <= saw_rom(399);
     when "000110010000" => data <= saw_rom(400);
     when "000110010001" => data <= saw_rom(401);
     when "000110010010" => data <= saw_rom(402);
     when "000110010011" => data <= saw_rom(403);
     when "000110010100" => data <= saw_rom(404);
     when "000110010101" => data <= saw_rom(405);
     when "000110010110" => data <= saw_rom(406);
     when "000110010111" => data <= saw_rom(407);
     when "000110011000" => data <= saw_rom(408);
     when "000110011001" => data <= saw_rom(409);
     when "000110011010" => data <= saw_rom(410);
     when "000110011011" => data <= saw_rom(411);
     when "000110011100" => data <= saw_rom(412);
     when "000110011101" => data <= saw_rom(413);
     when "000110011110" => data <= saw_rom(414);
     when "000110011111" => data <= saw_rom(415);
     when "000110100000" => data <= saw_rom(416);
     when "000110100001" => data <= saw_rom(417);
     when "000110100010" => data <= saw_rom(418);
     when "000110100011" => data <= saw_rom(419);
     when "000110100100" => data <= saw_rom(420);
     when "000110100101" => data <= saw_rom(421);
     when "000110100110" => data <= saw_rom(422);
     when "000110100111" => data <= saw_rom(423);
     when "000110101000" => data <= saw_rom(424);
     when "000110101001" => data <= saw_rom(425);
     when "000110101010" => data <= saw_rom(426);
     when "000110101011" => data <= saw_rom(427);
     when "000110101100" => data <= saw_rom(428);
     when "000110101101" => data <= saw_rom(429);
     when "000110101110" => data <= saw_rom(430);
     when "000110101111" => data <= saw_rom(431);
     when "000110110000" => data <= saw_rom(432);
     when "000110110001" => data <= saw_rom(433);
     when "000110110010" => data <= saw_rom(434);
     when "000110110011" => data <= saw_rom(435);
     when "000110110100" => data <= saw_rom(436);
     when "000110110101" => data <= saw_rom(437);
     when "000110110110" => data <= saw_rom(438);
     when "000110110111" => data <= saw_rom(439);
     when "000110111000" => data <= saw_rom(440);
     when "000110111001" => data <= saw_rom(441);
     when "000110111010" => data <= saw_rom(442);
     when "000110111011" => data <= saw_rom(443);
     when "000110111100" => data <= saw_rom(444);
     when "000110111101" => data <= saw_rom(445);
     when "000110111110" => data <= saw_rom(446);
     when "000110111111" => data <= saw_rom(447);
     when "000111000000" => data <= saw_rom(448);
     when "000111000001" => data <= saw_rom(449);
     when "000111000010" => data <= saw_rom(450);
     when "000111000011" => data <= saw_rom(451);
     when "000111000100" => data <= saw_rom(452);
     when "000111000101" => data <= saw_rom(453);
     when "000111000110" => data <= saw_rom(454);
     when "000111000111" => data <= saw_rom(455);
     when "000111001000" => data <= saw_rom(456);
     when "000111001001" => data <= saw_rom(457);
     when "000111001010" => data <= saw_rom(458);
     when "000111001011" => data <= saw_rom(459);
     when "000111001100" => data <= saw_rom(460);
     when "000111001101" => data <= saw_rom(461);
     when "000111001110" => data <= saw_rom(462);
     when "000111001111" => data <= saw_rom(463);
     when "000111010000" => data <= saw_rom(464);
     when "000111010001" => data <= saw_rom(465);
     when "000111010010" => data <= saw_rom(466);
     when "000111010011" => data <= saw_rom(467);
     when "000111010100" => data <= saw_rom(468);
     when "000111010101" => data <= saw_rom(469);
     when "000111010110" => data <= saw_rom(470);
     when "000111010111" => data <= saw_rom(471);
     when "000111011000" => data <= saw_rom(472);
     when "000111011001" => data <= saw_rom(473);
     when "000111011010" => data <= saw_rom(474);
     when "000111011011" => data <= saw_rom(475);
     when "000111011100" => data <= saw_rom(476);
     when "000111011101" => data <= saw_rom(477);
     when "000111011110" => data <= saw_rom(478);
     when "000111011111" => data <= saw_rom(479);
     when "000111100000" => data <= saw_rom(480);
     when "000111100001" => data <= saw_rom(481);
     when "000111100010" => data <= saw_rom(482);
     when "000111100011" => data <= saw_rom(483);
     when "000111100100" => data <= saw_rom(484);
     when "000111100101" => data <= saw_rom(485);
     when "000111100110" => data <= saw_rom(486);
     when "000111100111" => data <= saw_rom(487);
     when "000111101000" => data <= saw_rom(488);
     when "000111101001" => data <= saw_rom(489);
     when "000111101010" => data <= saw_rom(490);
     when "000111101011" => data <= saw_rom(491);
     when "000111101100" => data <= saw_rom(492);
     when "000111101101" => data <= saw_rom(493);
     when "000111101110" => data <= saw_rom(494);
     when "000111101111" => data <= saw_rom(495);
     when "000111110000" => data <= saw_rom(496);
     when "000111110001" => data <= saw_rom(497);
     when "000111110010" => data <= saw_rom(498);
     when "000111110011" => data <= saw_rom(499);
     when "000111110100" => data <= saw_rom(500);
     when "000111110101" => data <= saw_rom(501);
     when "000111110110" => data <= saw_rom(502);
     when "000111110111" => data <= saw_rom(503);
     when "000111111000" => data <= saw_rom(504);
     when "000111111001" => data <= saw_rom(505);
     when "000111111010" => data <= saw_rom(506);
     when "000111111011" => data <= saw_rom(507);
     when "000111111100" => data <= saw_rom(508);
     when "000111111101" => data <= saw_rom(509);
     when "000111111110" => data <= saw_rom(510);
     when "000111111111" => data <= saw_rom(511);
     when "001000000000" => data <= saw_rom(512);
     when "001000000001" => data <= saw_rom(513);
     when "001000000010" => data <= saw_rom(514);
     when "001000000011" => data <= saw_rom(515);
     when "001000000100" => data <= saw_rom(516);
     when "001000000101" => data <= saw_rom(517);
     when "001000000110" => data <= saw_rom(518);
     when "001000000111" => data <= saw_rom(519);
     when "001000001000" => data <= saw_rom(520);
     when "001000001001" => data <= saw_rom(521);
     when "001000001010" => data <= saw_rom(522);
     when "001000001011" => data <= saw_rom(523);
     when "001000001100" => data <= saw_rom(524);
     when "001000001101" => data <= saw_rom(525);
     when "001000001110" => data <= saw_rom(526);
     when "001000001111" => data <= saw_rom(527);
     when "001000010000" => data <= saw_rom(528);
     when "001000010001" => data <= saw_rom(529);
     when "001000010010" => data <= saw_rom(530);
     when "001000010011" => data <= saw_rom(531);
     when "001000010100" => data <= saw_rom(532);
     when "001000010101" => data <= saw_rom(533);
     when "001000010110" => data <= saw_rom(534);
     when "001000010111" => data <= saw_rom(535);
     when "001000011000" => data <= saw_rom(536);
     when "001000011001" => data <= saw_rom(537);
     when "001000011010" => data <= saw_rom(538);
     when "001000011011" => data <= saw_rom(539);
     when "001000011100" => data <= saw_rom(540);
     when "001000011101" => data <= saw_rom(541);
     when "001000011110" => data <= saw_rom(542);
     when "001000011111" => data <= saw_rom(543);
     when "001000100000" => data <= saw_rom(544);
     when "001000100001" => data <= saw_rom(545);
     when "001000100010" => data <= saw_rom(546);
     when "001000100011" => data <= saw_rom(547);
     when "001000100100" => data <= saw_rom(548);
     when "001000100101" => data <= saw_rom(549);
     when "001000100110" => data <= saw_rom(550);
     when "001000100111" => data <= saw_rom(551);
     when "001000101000" => data <= saw_rom(552);
     when "001000101001" => data <= saw_rom(553);
     when "001000101010" => data <= saw_rom(554);
     when "001000101011" => data <= saw_rom(555);
     when "001000101100" => data <= saw_rom(556);
     when "001000101101" => data <= saw_rom(557);
     when "001000101110" => data <= saw_rom(558);
     when "001000101111" => data <= saw_rom(559);
     when "001000110000" => data <= saw_rom(560);
     when "001000110001" => data <= saw_rom(561);
     when "001000110010" => data <= saw_rom(562);
     when "001000110011" => data <= saw_rom(563);
     when "001000110100" => data <= saw_rom(564);
     when "001000110101" => data <= saw_rom(565);
     when "001000110110" => data <= saw_rom(566);
     when "001000110111" => data <= saw_rom(567);
     when "001000111000" => data <= saw_rom(568);
     when "001000111001" => data <= saw_rom(569);
     when "001000111010" => data <= saw_rom(570);
     when "001000111011" => data <= saw_rom(571);
     when "001000111100" => data <= saw_rom(572);
     when "001000111101" => data <= saw_rom(573);
     when "001000111110" => data <= saw_rom(574);
     when "001000111111" => data <= saw_rom(575);
     when "001001000000" => data <= saw_rom(576);
     when "001001000001" => data <= saw_rom(577);
     when "001001000010" => data <= saw_rom(578);
     when "001001000011" => data <= saw_rom(579);
     when "001001000100" => data <= saw_rom(580);
     when "001001000101" => data <= saw_rom(581);
     when "001001000110" => data <= saw_rom(582);
     when "001001000111" => data <= saw_rom(583);
     when "001001001000" => data <= saw_rom(584);
     when "001001001001" => data <= saw_rom(585);
     when "001001001010" => data <= saw_rom(586);
     when "001001001011" => data <= saw_rom(587);
     when "001001001100" => data <= saw_rom(588);
     when "001001001101" => data <= saw_rom(589);
     when "001001001110" => data <= saw_rom(590);
     when "001001001111" => data <= saw_rom(591);
     when "001001010000" => data <= saw_rom(592);
     when "001001010001" => data <= saw_rom(593);
     when "001001010010" => data <= saw_rom(594);
     when "001001010011" => data <= saw_rom(595);
     when "001001010100" => data <= saw_rom(596);
     when "001001010101" => data <= saw_rom(597);
     when "001001010110" => data <= saw_rom(598);
     when "001001010111" => data <= saw_rom(599);
     when "001001011000" => data <= saw_rom(600);
     when "001001011001" => data <= saw_rom(601);
     when "001001011010" => data <= saw_rom(602);
     when "001001011011" => data <= saw_rom(603);
     when "001001011100" => data <= saw_rom(604);
     when "001001011101" => data <= saw_rom(605);
     when "001001011110" => data <= saw_rom(606);
     when "001001011111" => data <= saw_rom(607);
     when "001001100000" => data <= saw_rom(608);
     when "001001100001" => data <= saw_rom(609);
     when "001001100010" => data <= saw_rom(610);
     when "001001100011" => data <= saw_rom(611);
     when "001001100100" => data <= saw_rom(612);
     when "001001100101" => data <= saw_rom(613);
     when "001001100110" => data <= saw_rom(614);
     when "001001100111" => data <= saw_rom(615);
     when "001001101000" => data <= saw_rom(616);
     when "001001101001" => data <= saw_rom(617);
     when "001001101010" => data <= saw_rom(618);
     when "001001101011" => data <= saw_rom(619);
     when "001001101100" => data <= saw_rom(620);
     when "001001101101" => data <= saw_rom(621);
     when "001001101110" => data <= saw_rom(622);
     when "001001101111" => data <= saw_rom(623);
     when "001001110000" => data <= saw_rom(624);
     when "001001110001" => data <= saw_rom(625);
     when "001001110010" => data <= saw_rom(626);
     when "001001110011" => data <= saw_rom(627);
     when "001001110100" => data <= saw_rom(628);
     when "001001110101" => data <= saw_rom(629);
     when "001001110110" => data <= saw_rom(630);
     when "001001110111" => data <= saw_rom(631);
     when "001001111000" => data <= saw_rom(632);
     when "001001111001" => data <= saw_rom(633);
     when "001001111010" => data <= saw_rom(634);
     when "001001111011" => data <= saw_rom(635);
     when "001001111100" => data <= saw_rom(636);
     when "001001111101" => data <= saw_rom(637);
     when "001001111110" => data <= saw_rom(638);
     when "001001111111" => data <= saw_rom(639);
     when "001010000000" => data <= saw_rom(640);
     when "001010000001" => data <= saw_rom(641);
     when "001010000010" => data <= saw_rom(642);
     when "001010000011" => data <= saw_rom(643);
     when "001010000100" => data <= saw_rom(644);
     when "001010000101" => data <= saw_rom(645);
     when "001010000110" => data <= saw_rom(646);
     when "001010000111" => data <= saw_rom(647);
     when "001010001000" => data <= saw_rom(648);
     when "001010001001" => data <= saw_rom(649);
     when "001010001010" => data <= saw_rom(650);
     when "001010001011" => data <= saw_rom(651);
     when "001010001100" => data <= saw_rom(652);
     when "001010001101" => data <= saw_rom(653);
     when "001010001110" => data <= saw_rom(654);
     when "001010001111" => data <= saw_rom(655);
     when "001010010000" => data <= saw_rom(656);
     when "001010010001" => data <= saw_rom(657);
     when "001010010010" => data <= saw_rom(658);
     when "001010010011" => data <= saw_rom(659);
     when "001010010100" => data <= saw_rom(660);
     when "001010010101" => data <= saw_rom(661);
     when "001010010110" => data <= saw_rom(662);
     when "001010010111" => data <= saw_rom(663);
     when "001010011000" => data <= saw_rom(664);
     when "001010011001" => data <= saw_rom(665);
     when "001010011010" => data <= saw_rom(666);
     when "001010011011" => data <= saw_rom(667);
     when "001010011100" => data <= saw_rom(668);
     when "001010011101" => data <= saw_rom(669);
     when "001010011110" => data <= saw_rom(670);
     when "001010011111" => data <= saw_rom(671);
     when "001010100000" => data <= saw_rom(672);
     when "001010100001" => data <= saw_rom(673);
     when "001010100010" => data <= saw_rom(674);
     when "001010100011" => data <= saw_rom(675);
     when "001010100100" => data <= saw_rom(676);
     when "001010100101" => data <= saw_rom(677);
     when "001010100110" => data <= saw_rom(678);
     when "001010100111" => data <= saw_rom(679);
     when "001010101000" => data <= saw_rom(680);
     when "001010101001" => data <= saw_rom(681);
     when "001010101010" => data <= saw_rom(682);
     when "001010101011" => data <= saw_rom(683);
     when "001010101100" => data <= saw_rom(684);
     when "001010101101" => data <= saw_rom(685);
     when "001010101110" => data <= saw_rom(686);
     when "001010101111" => data <= saw_rom(687);
     when "001010110000" => data <= saw_rom(688);
     when "001010110001" => data <= saw_rom(689);
     when "001010110010" => data <= saw_rom(690);
     when "001010110011" => data <= saw_rom(691);
     when "001010110100" => data <= saw_rom(692);
     when "001010110101" => data <= saw_rom(693);
     when "001010110110" => data <= saw_rom(694);
     when "001010110111" => data <= saw_rom(695);
     when "001010111000" => data <= saw_rom(696);
     when "001010111001" => data <= saw_rom(697);
     when "001010111010" => data <= saw_rom(698);
     when "001010111011" => data <= saw_rom(699);
     when "001010111100" => data <= saw_rom(700);
     when "001010111101" => data <= saw_rom(701);
     when "001010111110" => data <= saw_rom(702);
     when "001010111111" => data <= saw_rom(703);
     when "001011000000" => data <= saw_rom(704);
     when "001011000001" => data <= saw_rom(705);
     when "001011000010" => data <= saw_rom(706);
     when "001011000011" => data <= saw_rom(707);
     when "001011000100" => data <= saw_rom(708);
     when "001011000101" => data <= saw_rom(709);
     when "001011000110" => data <= saw_rom(710);
     when "001011000111" => data <= saw_rom(711);
     when "001011001000" => data <= saw_rom(712);
     when "001011001001" => data <= saw_rom(713);
     when "001011001010" => data <= saw_rom(714);
     when "001011001011" => data <= saw_rom(715);
     when "001011001100" => data <= saw_rom(716);
     when "001011001101" => data <= saw_rom(717);
     when "001011001110" => data <= saw_rom(718);
     when "001011001111" => data <= saw_rom(719);
     when "001011010000" => data <= saw_rom(720);
     when "001011010001" => data <= saw_rom(721);
     when "001011010010" => data <= saw_rom(722);
     when "001011010011" => data <= saw_rom(723);
     when "001011010100" => data <= saw_rom(724);
     when "001011010101" => data <= saw_rom(725);
     when "001011010110" => data <= saw_rom(726);
     when "001011010111" => data <= saw_rom(727);
     when "001011011000" => data <= saw_rom(728);
     when "001011011001" => data <= saw_rom(729);
     when "001011011010" => data <= saw_rom(730);
     when "001011011011" => data <= saw_rom(731);
     when "001011011100" => data <= saw_rom(732);
     when "001011011101" => data <= saw_rom(733);
     when "001011011110" => data <= saw_rom(734);
     when "001011011111" => data <= saw_rom(735);
     when "001011100000" => data <= saw_rom(736);
     when "001011100001" => data <= saw_rom(737);
     when "001011100010" => data <= saw_rom(738);
     when "001011100011" => data <= saw_rom(739);
     when "001011100100" => data <= saw_rom(740);
     when "001011100101" => data <= saw_rom(741);
     when "001011100110" => data <= saw_rom(742);
     when "001011100111" => data <= saw_rom(743);
     when "001011101000" => data <= saw_rom(744);
     when "001011101001" => data <= saw_rom(745);
     when "001011101010" => data <= saw_rom(746);
     when "001011101011" => data <= saw_rom(747);
     when "001011101100" => data <= saw_rom(748);
     when "001011101101" => data <= saw_rom(749);
     when "001011101110" => data <= saw_rom(750);
     when "001011101111" => data <= saw_rom(751);
     when "001011110000" => data <= saw_rom(752);
     when "001011110001" => data <= saw_rom(753);
     when "001011110010" => data <= saw_rom(754);
     when "001011110011" => data <= saw_rom(755);
     when "001011110100" => data <= saw_rom(756);
     when "001011110101" => data <= saw_rom(757);
     when "001011110110" => data <= saw_rom(758);
     when "001011110111" => data <= saw_rom(759);
     when "001011111000" => data <= saw_rom(760);
     when "001011111001" => data <= saw_rom(761);
     when "001011111010" => data <= saw_rom(762);
     when "001011111011" => data <= saw_rom(763);
     when "001011111100" => data <= saw_rom(764);
     when "001011111101" => data <= saw_rom(765);
     when "001011111110" => data <= saw_rom(766);
     when "001011111111" => data <= saw_rom(767);
     when "001100000000" => data <= saw_rom(768);
     when "001100000001" => data <= saw_rom(769);
     when "001100000010" => data <= saw_rom(770);
     when "001100000011" => data <= saw_rom(771);
     when "001100000100" => data <= saw_rom(772);
     when "001100000101" => data <= saw_rom(773);
     when "001100000110" => data <= saw_rom(774);
     when "001100000111" => data <= saw_rom(775);
     when "001100001000" => data <= saw_rom(776);
     when "001100001001" => data <= saw_rom(777);
     when "001100001010" => data <= saw_rom(778);
     when "001100001011" => data <= saw_rom(779);
     when "001100001100" => data <= saw_rom(780);
     when "001100001101" => data <= saw_rom(781);
     when "001100001110" => data <= saw_rom(782);
     when "001100001111" => data <= saw_rom(783);
     when "001100010000" => data <= saw_rom(784);
     when "001100010001" => data <= saw_rom(785);
     when "001100010010" => data <= saw_rom(786);
     when "001100010011" => data <= saw_rom(787);
     when "001100010100" => data <= saw_rom(788);
     when "001100010101" => data <= saw_rom(789);
     when "001100010110" => data <= saw_rom(790);
     when "001100010111" => data <= saw_rom(791);
     when "001100011000" => data <= saw_rom(792);
     when "001100011001" => data <= saw_rom(793);
     when "001100011010" => data <= saw_rom(794);
     when "001100011011" => data <= saw_rom(795);
     when "001100011100" => data <= saw_rom(796);
     when "001100011101" => data <= saw_rom(797);
     when "001100011110" => data <= saw_rom(798);
     when "001100011111" => data <= saw_rom(799);
     when "001100100000" => data <= saw_rom(800);
     when "001100100001" => data <= saw_rom(801);
     when "001100100010" => data <= saw_rom(802);
     when "001100100011" => data <= saw_rom(803);
     when "001100100100" => data <= saw_rom(804);
     when "001100100101" => data <= saw_rom(805);
     when "001100100110" => data <= saw_rom(806);
     when "001100100111" => data <= saw_rom(807);
     when "001100101000" => data <= saw_rom(808);
     when "001100101001" => data <= saw_rom(809);
     when "001100101010" => data <= saw_rom(810);
     when "001100101011" => data <= saw_rom(811);
     when "001100101100" => data <= saw_rom(812);
     when "001100101101" => data <= saw_rom(813);
     when "001100101110" => data <= saw_rom(814);
     when "001100101111" => data <= saw_rom(815);
     when "001100110000" => data <= saw_rom(816);
     when "001100110001" => data <= saw_rom(817);
     when "001100110010" => data <= saw_rom(818);
     when "001100110011" => data <= saw_rom(819);
     when "001100110100" => data <= saw_rom(820);
     when "001100110101" => data <= saw_rom(821);
     when "001100110110" => data <= saw_rom(822);
     when "001100110111" => data <= saw_rom(823);
     when "001100111000" => data <= saw_rom(824);
     when "001100111001" => data <= saw_rom(825);
     when "001100111010" => data <= saw_rom(826);
     when "001100111011" => data <= saw_rom(827);
     when "001100111100" => data <= saw_rom(828);
     when "001100111101" => data <= saw_rom(829);
     when "001100111110" => data <= saw_rom(830);
     when "001100111111" => data <= saw_rom(831);
     when "001101000000" => data <= saw_rom(832);
     when "001101000001" => data <= saw_rom(833);
     when "001101000010" => data <= saw_rom(834);
     when "001101000011" => data <= saw_rom(835);
     when "001101000100" => data <= saw_rom(836);
     when "001101000101" => data <= saw_rom(837);
     when "001101000110" => data <= saw_rom(838);
     when "001101000111" => data <= saw_rom(839);
     when "001101001000" => data <= saw_rom(840);
     when "001101001001" => data <= saw_rom(841);
     when "001101001010" => data <= saw_rom(842);
     when "001101001011" => data <= saw_rom(843);
     when "001101001100" => data <= saw_rom(844);
     when "001101001101" => data <= saw_rom(845);
     when "001101001110" => data <= saw_rom(846);
     when "001101001111" => data <= saw_rom(847);
     when "001101010000" => data <= saw_rom(848);
     when "001101010001" => data <= saw_rom(849);
     when "001101010010" => data <= saw_rom(850);
     when "001101010011" => data <= saw_rom(851);
     when "001101010100" => data <= saw_rom(852);
     when "001101010101" => data <= saw_rom(853);
     when "001101010110" => data <= saw_rom(854);
     when "001101010111" => data <= saw_rom(855);
     when "001101011000" => data <= saw_rom(856);
     when "001101011001" => data <= saw_rom(857);
     when "001101011010" => data <= saw_rom(858);
     when "001101011011" => data <= saw_rom(859);
     when "001101011100" => data <= saw_rom(860);
     when "001101011101" => data <= saw_rom(861);
     when "001101011110" => data <= saw_rom(862);
     when "001101011111" => data <= saw_rom(863);
     when "001101100000" => data <= saw_rom(864);
     when "001101100001" => data <= saw_rom(865);
     when "001101100010" => data <= saw_rom(866);
     when "001101100011" => data <= saw_rom(867);
     when "001101100100" => data <= saw_rom(868);
     when "001101100101" => data <= saw_rom(869);
     when "001101100110" => data <= saw_rom(870);
     when "001101100111" => data <= saw_rom(871);
     when "001101101000" => data <= saw_rom(872);
     when "001101101001" => data <= saw_rom(873);
     when "001101101010" => data <= saw_rom(874);
     when "001101101011" => data <= saw_rom(875);
     when "001101101100" => data <= saw_rom(876);
     when "001101101101" => data <= saw_rom(877);
     when "001101101110" => data <= saw_rom(878);
     when "001101101111" => data <= saw_rom(879);
     when "001101110000" => data <= saw_rom(880);
     when "001101110001" => data <= saw_rom(881);
     when "001101110010" => data <= saw_rom(882);
     when "001101110011" => data <= saw_rom(883);
     when "001101110100" => data <= saw_rom(884);
     when "001101110101" => data <= saw_rom(885);
     when "001101110110" => data <= saw_rom(886);
     when "001101110111" => data <= saw_rom(887);
     when "001101111000" => data <= saw_rom(888);
     when "001101111001" => data <= saw_rom(889);
     when "001101111010" => data <= saw_rom(890);
     when "001101111011" => data <= saw_rom(891);
     when "001101111100" => data <= saw_rom(892);
     when "001101111101" => data <= saw_rom(893);
     when "001101111110" => data <= saw_rom(894);
     when "001101111111" => data <= saw_rom(895);
     when "001110000000" => data <= saw_rom(896);
     when "001110000001" => data <= saw_rom(897);
     when "001110000010" => data <= saw_rom(898);
     when "001110000011" => data <= saw_rom(899);
     when "001110000100" => data <= saw_rom(900);
     when "001110000101" => data <= saw_rom(901);
     when "001110000110" => data <= saw_rom(902);
     when "001110000111" => data <= saw_rom(903);
     when "001110001000" => data <= saw_rom(904);
     when "001110001001" => data <= saw_rom(905);
     when "001110001010" => data <= saw_rom(906);
     when "001110001011" => data <= saw_rom(907);
     when "001110001100" => data <= saw_rom(908);
     when "001110001101" => data <= saw_rom(909);
     when "001110001110" => data <= saw_rom(910);
     when "001110001111" => data <= saw_rom(911);
     when "001110010000" => data <= saw_rom(912);
     when "001110010001" => data <= saw_rom(913);
     when "001110010010" => data <= saw_rom(914);
     when "001110010011" => data <= saw_rom(915);
     when "001110010100" => data <= saw_rom(916);
     when "001110010101" => data <= saw_rom(917);
     when "001110010110" => data <= saw_rom(918);
     when "001110010111" => data <= saw_rom(919);
     when "001110011000" => data <= saw_rom(920);
     when "001110011001" => data <= saw_rom(921);
     when "001110011010" => data <= saw_rom(922);
     when "001110011011" => data <= saw_rom(923);
     when "001110011100" => data <= saw_rom(924);
     when "001110011101" => data <= saw_rom(925);
     when "001110011110" => data <= saw_rom(926);
     when "001110011111" => data <= saw_rom(927);
     when "001110100000" => data <= saw_rom(928);
     when "001110100001" => data <= saw_rom(929);
     when "001110100010" => data <= saw_rom(930);
     when "001110100011" => data <= saw_rom(931);
     when "001110100100" => data <= saw_rom(932);
     when "001110100101" => data <= saw_rom(933);
     when "001110100110" => data <= saw_rom(934);
     when "001110100111" => data <= saw_rom(935);
     when "001110101000" => data <= saw_rom(936);
     when "001110101001" => data <= saw_rom(937);
     when "001110101010" => data <= saw_rom(938);
     when "001110101011" => data <= saw_rom(939);
     when "001110101100" => data <= saw_rom(940);
     when "001110101101" => data <= saw_rom(941);
     when "001110101110" => data <= saw_rom(942);
     when "001110101111" => data <= saw_rom(943);
     when "001110110000" => data <= saw_rom(944);
     when "001110110001" => data <= saw_rom(945);
     when "001110110010" => data <= saw_rom(946);
     when "001110110011" => data <= saw_rom(947);
     when "001110110100" => data <= saw_rom(948);
     when "001110110101" => data <= saw_rom(949);
     when "001110110110" => data <= saw_rom(950);
     when "001110110111" => data <= saw_rom(951);
     when "001110111000" => data <= saw_rom(952);
     when "001110111001" => data <= saw_rom(953);
     when "001110111010" => data <= saw_rom(954);
     when "001110111011" => data <= saw_rom(955);
     when "001110111100" => data <= saw_rom(956);
     when "001110111101" => data <= saw_rom(957);
     when "001110111110" => data <= saw_rom(958);
     when "001110111111" => data <= saw_rom(959);
     when "001111000000" => data <= saw_rom(960);
     when "001111000001" => data <= saw_rom(961);
     when "001111000010" => data <= saw_rom(962);
     when "001111000011" => data <= saw_rom(963);
     when "001111000100" => data <= saw_rom(964);
     when "001111000101" => data <= saw_rom(965);
     when "001111000110" => data <= saw_rom(966);
     when "001111000111" => data <= saw_rom(967);
     when "001111001000" => data <= saw_rom(968);
     when "001111001001" => data <= saw_rom(969);
     when "001111001010" => data <= saw_rom(970);
     when "001111001011" => data <= saw_rom(971);
     when "001111001100" => data <= saw_rom(972);
     when "001111001101" => data <= saw_rom(973);
     when "001111001110" => data <= saw_rom(974);
     when "001111001111" => data <= saw_rom(975);
     when "001111010000" => data <= saw_rom(976);
     when "001111010001" => data <= saw_rom(977);
     when "001111010010" => data <= saw_rom(978);
     when "001111010011" => data <= saw_rom(979);
     when "001111010100" => data <= saw_rom(980);
     when "001111010101" => data <= saw_rom(981);
     when "001111010110" => data <= saw_rom(982);
     when "001111010111" => data <= saw_rom(983);
     when "001111011000" => data <= saw_rom(984);
     when "001111011001" => data <= saw_rom(985);
     when "001111011010" => data <= saw_rom(986);
     when "001111011011" => data <= saw_rom(987);
     when "001111011100" => data <= saw_rom(988);
     when "001111011101" => data <= saw_rom(989);
     when "001111011110" => data <= saw_rom(990);
     when "001111011111" => data <= saw_rom(991);
     when "001111100000" => data <= saw_rom(992);
     when "001111100001" => data <= saw_rom(993);
     when "001111100010" => data <= saw_rom(994);
     when "001111100011" => data <= saw_rom(995);
     when "001111100100" => data <= saw_rom(996);
     when "001111100101" => data <= saw_rom(997);
     when "001111100110" => data <= saw_rom(998);
     when "001111100111" => data <= saw_rom(999);
     when "001111101000" => data <= saw_rom(1000);
     when "001111101001" => data <= saw_rom(1001);
     when "001111101010" => data <= saw_rom(1002);
     when "001111101011" => data <= saw_rom(1003);
     when "001111101100" => data <= saw_rom(1004);
     when "001111101101" => data <= saw_rom(1005);
     when "001111101110" => data <= saw_rom(1006);
     when "001111101111" => data <= saw_rom(1007);
     when "001111110000" => data <= saw_rom(1008);
     when "001111110001" => data <= saw_rom(1009);
     when "001111110010" => data <= saw_rom(1010);
     when "001111110011" => data <= saw_rom(1011);
     when "001111110100" => data <= saw_rom(1012);
     when "001111110101" => data <= saw_rom(1013);
     when "001111110110" => data <= saw_rom(1014);
     when "001111110111" => data <= saw_rom(1015);
     when "001111111000" => data <= saw_rom(1016);
     when "001111111001" => data <= saw_rom(1017);
     when "001111111010" => data <= saw_rom(1018);
     when "001111111011" => data <= saw_rom(1019);
     when "001111111100" => data <= saw_rom(1020);
     when "001111111101" => data <= saw_rom(1021);
     when "001111111110" => data <= saw_rom(1022);
     when "001111111111" => data <= saw_rom(1023);
     when "010000000000" => data <= saw_rom(1024);
     when "010000000001" => data <= saw_rom(1025);
     when "010000000010" => data <= saw_rom(1026);
     when "010000000011" => data <= saw_rom(1027);
     when "010000000100" => data <= saw_rom(1028);
     when "010000000101" => data <= saw_rom(1029);
     when "010000000110" => data <= saw_rom(1030);
     when "010000000111" => data <= saw_rom(1031);
     when "010000001000" => data <= saw_rom(1032);
     when "010000001001" => data <= saw_rom(1033);
     when "010000001010" => data <= saw_rom(1034);
     when "010000001011" => data <= saw_rom(1035);
     when "010000001100" => data <= saw_rom(1036);
     when "010000001101" => data <= saw_rom(1037);
     when "010000001110" => data <= saw_rom(1038);
     when "010000001111" => data <= saw_rom(1039);
     when "010000010000" => data <= saw_rom(1040);
     when "010000010001" => data <= saw_rom(1041);
     when "010000010010" => data <= saw_rom(1042);
     when "010000010011" => data <= saw_rom(1043);
     when "010000010100" => data <= saw_rom(1044);
     when "010000010101" => data <= saw_rom(1045);
     when "010000010110" => data <= saw_rom(1046);
     when "010000010111" => data <= saw_rom(1047);
     when "010000011000" => data <= saw_rom(1048);
     when "010000011001" => data <= saw_rom(1049);
     when "010000011010" => data <= saw_rom(1050);
     when "010000011011" => data <= saw_rom(1051);
     when "010000011100" => data <= saw_rom(1052);
     when "010000011101" => data <= saw_rom(1053);
     when "010000011110" => data <= saw_rom(1054);
     when "010000011111" => data <= saw_rom(1055);
     when "010000100000" => data <= saw_rom(1056);
     when "010000100001" => data <= saw_rom(1057);
     when "010000100010" => data <= saw_rom(1058);
     when "010000100011" => data <= saw_rom(1059);
     when "010000100100" => data <= saw_rom(1060);
     when "010000100101" => data <= saw_rom(1061);
     when "010000100110" => data <= saw_rom(1062);
     when "010000100111" => data <= saw_rom(1063);
     when "010000101000" => data <= saw_rom(1064);
     when "010000101001" => data <= saw_rom(1065);
     when "010000101010" => data <= saw_rom(1066);
     when "010000101011" => data <= saw_rom(1067);
     when "010000101100" => data <= saw_rom(1068);
     when "010000101101" => data <= saw_rom(1069);
     when "010000101110" => data <= saw_rom(1070);
     when "010000101111" => data <= saw_rom(1071);
     when "010000110000" => data <= saw_rom(1072);
     when "010000110001" => data <= saw_rom(1073);
     when "010000110010" => data <= saw_rom(1074);
     when "010000110011" => data <= saw_rom(1075);
     when "010000110100" => data <= saw_rom(1076);
     when "010000110101" => data <= saw_rom(1077);
     when "010000110110" => data <= saw_rom(1078);
     when "010000110111" => data <= saw_rom(1079);
     when "010000111000" => data <= saw_rom(1080);
     when "010000111001" => data <= saw_rom(1081);
     when "010000111010" => data <= saw_rom(1082);
     when "010000111011" => data <= saw_rom(1083);
     when "010000111100" => data <= saw_rom(1084);
     when "010000111101" => data <= saw_rom(1085);
     when "010000111110" => data <= saw_rom(1086);
     when "010000111111" => data <= saw_rom(1087);
     when "010001000000" => data <= saw_rom(1088);
     when "010001000001" => data <= saw_rom(1089);
     when "010001000010" => data <= saw_rom(1090);
     when "010001000011" => data <= saw_rom(1091);
     when "010001000100" => data <= saw_rom(1092);
     when "010001000101" => data <= saw_rom(1093);
     when "010001000110" => data <= saw_rom(1094);
     when "010001000111" => data <= saw_rom(1095);
     when "010001001000" => data <= saw_rom(1096);
     when "010001001001" => data <= saw_rom(1097);
     when "010001001010" => data <= saw_rom(1098);
     when "010001001011" => data <= saw_rom(1099);
     when "010001001100" => data <= saw_rom(1100);
     when "010001001101" => data <= saw_rom(1101);
     when "010001001110" => data <= saw_rom(1102);
     when "010001001111" => data <= saw_rom(1103);
     when "010001010000" => data <= saw_rom(1104);
     when "010001010001" => data <= saw_rom(1105);
     when "010001010010" => data <= saw_rom(1106);
     when "010001010011" => data <= saw_rom(1107);
     when "010001010100" => data <= saw_rom(1108);
     when "010001010101" => data <= saw_rom(1109);
     when "010001010110" => data <= saw_rom(1110);
     when "010001010111" => data <= saw_rom(1111);
     when "010001011000" => data <= saw_rom(1112);
     when "010001011001" => data <= saw_rom(1113);
     when "010001011010" => data <= saw_rom(1114);
     when "010001011011" => data <= saw_rom(1115);
     when "010001011100" => data <= saw_rom(1116);
     when "010001011101" => data <= saw_rom(1117);
     when "010001011110" => data <= saw_rom(1118);
     when "010001011111" => data <= saw_rom(1119);
     when "010001100000" => data <= saw_rom(1120);
     when "010001100001" => data <= saw_rom(1121);
     when "010001100010" => data <= saw_rom(1122);
     when "010001100011" => data <= saw_rom(1123);
     when "010001100100" => data <= saw_rom(1124);
     when "010001100101" => data <= saw_rom(1125);
     when "010001100110" => data <= saw_rom(1126);
     when "010001100111" => data <= saw_rom(1127);
     when "010001101000" => data <= saw_rom(1128);
     when "010001101001" => data <= saw_rom(1129);
     when "010001101010" => data <= saw_rom(1130);
     when "010001101011" => data <= saw_rom(1131);
     when "010001101100" => data <= saw_rom(1132);
     when "010001101101" => data <= saw_rom(1133);
     when "010001101110" => data <= saw_rom(1134);
     when "010001101111" => data <= saw_rom(1135);
     when "010001110000" => data <= saw_rom(1136);
     when "010001110001" => data <= saw_rom(1137);
     when "010001110010" => data <= saw_rom(1138);
     when "010001110011" => data <= saw_rom(1139);
     when "010001110100" => data <= saw_rom(1140);
     when "010001110101" => data <= saw_rom(1141);
     when "010001110110" => data <= saw_rom(1142);
     when "010001110111" => data <= saw_rom(1143);
     when "010001111000" => data <= saw_rom(1144);
     when "010001111001" => data <= saw_rom(1145);
     when "010001111010" => data <= saw_rom(1146);
     when "010001111011" => data <= saw_rom(1147);
     when "010001111100" => data <= saw_rom(1148);
     when "010001111101" => data <= saw_rom(1149);
     when "010001111110" => data <= saw_rom(1150);
     when "010001111111" => data <= saw_rom(1151);
     when "010010000000" => data <= saw_rom(1152);
     when "010010000001" => data <= saw_rom(1153);
     when "010010000010" => data <= saw_rom(1154);
     when "010010000011" => data <= saw_rom(1155);
     when "010010000100" => data <= saw_rom(1156);
     when "010010000101" => data <= saw_rom(1157);
     when "010010000110" => data <= saw_rom(1158);
     when "010010000111" => data <= saw_rom(1159);
     when "010010001000" => data <= saw_rom(1160);
     when "010010001001" => data <= saw_rom(1161);
     when "010010001010" => data <= saw_rom(1162);
     when "010010001011" => data <= saw_rom(1163);
     when "010010001100" => data <= saw_rom(1164);
     when "010010001101" => data <= saw_rom(1165);
     when "010010001110" => data <= saw_rom(1166);
     when "010010001111" => data <= saw_rom(1167);
     when "010010010000" => data <= saw_rom(1168);
     when "010010010001" => data <= saw_rom(1169);
     when "010010010010" => data <= saw_rom(1170);
     when "010010010011" => data <= saw_rom(1171);
     when "010010010100" => data <= saw_rom(1172);
     when "010010010101" => data <= saw_rom(1173);
     when "010010010110" => data <= saw_rom(1174);
     when "010010010111" => data <= saw_rom(1175);
     when "010010011000" => data <= saw_rom(1176);
     when "010010011001" => data <= saw_rom(1177);
     when "010010011010" => data <= saw_rom(1178);
     when "010010011011" => data <= saw_rom(1179);
     when "010010011100" => data <= saw_rom(1180);
     when "010010011101" => data <= saw_rom(1181);
     when "010010011110" => data <= saw_rom(1182);
     when "010010011111" => data <= saw_rom(1183);
     when "010010100000" => data <= saw_rom(1184);
     when "010010100001" => data <= saw_rom(1185);
     when "010010100010" => data <= saw_rom(1186);
     when "010010100011" => data <= saw_rom(1187);
     when "010010100100" => data <= saw_rom(1188);
     when "010010100101" => data <= saw_rom(1189);
     when "010010100110" => data <= saw_rom(1190);
     when "010010100111" => data <= saw_rom(1191);
     when "010010101000" => data <= saw_rom(1192);
     when "010010101001" => data <= saw_rom(1193);
     when "010010101010" => data <= saw_rom(1194);
     when "010010101011" => data <= saw_rom(1195);
     when "010010101100" => data <= saw_rom(1196);
     when "010010101101" => data <= saw_rom(1197);
     when "010010101110" => data <= saw_rom(1198);
     when "010010101111" => data <= saw_rom(1199);
     when "010010110000" => data <= saw_rom(1200);
     when "010010110001" => data <= saw_rom(1201);
     when "010010110010" => data <= saw_rom(1202);
     when "010010110011" => data <= saw_rom(1203);
     when "010010110100" => data <= saw_rom(1204);
     when "010010110101" => data <= saw_rom(1205);
     when "010010110110" => data <= saw_rom(1206);
     when "010010110111" => data <= saw_rom(1207);
     when "010010111000" => data <= saw_rom(1208);
     when "010010111001" => data <= saw_rom(1209);
     when "010010111010" => data <= saw_rom(1210);
     when "010010111011" => data <= saw_rom(1211);
     when "010010111100" => data <= saw_rom(1212);
     when "010010111101" => data <= saw_rom(1213);
     when "010010111110" => data <= saw_rom(1214);
     when "010010111111" => data <= saw_rom(1215);
     when "010011000000" => data <= saw_rom(1216);
     when "010011000001" => data <= saw_rom(1217);
     when "010011000010" => data <= saw_rom(1218);
     when "010011000011" => data <= saw_rom(1219);
     when "010011000100" => data <= saw_rom(1220);
     when "010011000101" => data <= saw_rom(1221);
     when "010011000110" => data <= saw_rom(1222);
     when "010011000111" => data <= saw_rom(1223);
     when "010011001000" => data <= saw_rom(1224);
     when "010011001001" => data <= saw_rom(1225);
     when "010011001010" => data <= saw_rom(1226);
     when "010011001011" => data <= saw_rom(1227);
     when "010011001100" => data <= saw_rom(1228);
     when "010011001101" => data <= saw_rom(1229);
     when "010011001110" => data <= saw_rom(1230);
     when "010011001111" => data <= saw_rom(1231);
     when "010011010000" => data <= saw_rom(1232);
     when "010011010001" => data <= saw_rom(1233);
     when "010011010010" => data <= saw_rom(1234);
     when "010011010011" => data <= saw_rom(1235);
     when "010011010100" => data <= saw_rom(1236);
     when "010011010101" => data <= saw_rom(1237);
     when "010011010110" => data <= saw_rom(1238);
     when "010011010111" => data <= saw_rom(1239);
     when "010011011000" => data <= saw_rom(1240);
     when "010011011001" => data <= saw_rom(1241);
     when "010011011010" => data <= saw_rom(1242);
     when "010011011011" => data <= saw_rom(1243);
     when "010011011100" => data <= saw_rom(1244);
     when "010011011101" => data <= saw_rom(1245);
     when "010011011110" => data <= saw_rom(1246);
     when "010011011111" => data <= saw_rom(1247);
     when "010011100000" => data <= saw_rom(1248);
     when "010011100001" => data <= saw_rom(1249);
     when "010011100010" => data <= saw_rom(1250);
     when "010011100011" => data <= saw_rom(1251);
     when "010011100100" => data <= saw_rom(1252);
     when "010011100101" => data <= saw_rom(1253);
     when "010011100110" => data <= saw_rom(1254);
     when "010011100111" => data <= saw_rom(1255);
     when "010011101000" => data <= saw_rom(1256);
     when "010011101001" => data <= saw_rom(1257);
     when "010011101010" => data <= saw_rom(1258);
     when "010011101011" => data <= saw_rom(1259);
     when "010011101100" => data <= saw_rom(1260);
     when "010011101101" => data <= saw_rom(1261);
     when "010011101110" => data <= saw_rom(1262);
     when "010011101111" => data <= saw_rom(1263);
     when "010011110000" => data <= saw_rom(1264);
     when "010011110001" => data <= saw_rom(1265);
     when "010011110010" => data <= saw_rom(1266);
     when "010011110011" => data <= saw_rom(1267);
     when "010011110100" => data <= saw_rom(1268);
     when "010011110101" => data <= saw_rom(1269);
     when "010011110110" => data <= saw_rom(1270);
     when "010011110111" => data <= saw_rom(1271);
     when "010011111000" => data <= saw_rom(1272);
     when "010011111001" => data <= saw_rom(1273);
     when "010011111010" => data <= saw_rom(1274);
     when "010011111011" => data <= saw_rom(1275);
     when "010011111100" => data <= saw_rom(1276);
     when "010011111101" => data <= saw_rom(1277);
     when "010011111110" => data <= saw_rom(1278);
     when "010011111111" => data <= saw_rom(1279);
     when "010100000000" => data <= saw_rom(1280);
     when "010100000001" => data <= saw_rom(1281);
     when "010100000010" => data <= saw_rom(1282);
     when "010100000011" => data <= saw_rom(1283);
     when "010100000100" => data <= saw_rom(1284);
     when "010100000101" => data <= saw_rom(1285);
     when "010100000110" => data <= saw_rom(1286);
     when "010100000111" => data <= saw_rom(1287);
     when "010100001000" => data <= saw_rom(1288);
     when "010100001001" => data <= saw_rom(1289);
     when "010100001010" => data <= saw_rom(1290);
     when "010100001011" => data <= saw_rom(1291);
     when "010100001100" => data <= saw_rom(1292);
     when "010100001101" => data <= saw_rom(1293);
     when "010100001110" => data <= saw_rom(1294);
     when "010100001111" => data <= saw_rom(1295);
     when "010100010000" => data <= saw_rom(1296);
     when "010100010001" => data <= saw_rom(1297);
     when "010100010010" => data <= saw_rom(1298);
     when "010100010011" => data <= saw_rom(1299);
     when "010100010100" => data <= saw_rom(1300);
     when "010100010101" => data <= saw_rom(1301);
     when "010100010110" => data <= saw_rom(1302);
     when "010100010111" => data <= saw_rom(1303);
     when "010100011000" => data <= saw_rom(1304);
     when "010100011001" => data <= saw_rom(1305);
     when "010100011010" => data <= saw_rom(1306);
     when "010100011011" => data <= saw_rom(1307);
     when "010100011100" => data <= saw_rom(1308);
     when "010100011101" => data <= saw_rom(1309);
     when "010100011110" => data <= saw_rom(1310);
     when "010100011111" => data <= saw_rom(1311);
     when "010100100000" => data <= saw_rom(1312);
     when "010100100001" => data <= saw_rom(1313);
     when "010100100010" => data <= saw_rom(1314);
     when "010100100011" => data <= saw_rom(1315);
     when "010100100100" => data <= saw_rom(1316);
     when "010100100101" => data <= saw_rom(1317);
     when "010100100110" => data <= saw_rom(1318);
     when "010100100111" => data <= saw_rom(1319);
     when "010100101000" => data <= saw_rom(1320);
     when "010100101001" => data <= saw_rom(1321);
     when "010100101010" => data <= saw_rom(1322);
     when "010100101011" => data <= saw_rom(1323);
     when "010100101100" => data <= saw_rom(1324);
     when "010100101101" => data <= saw_rom(1325);
     when "010100101110" => data <= saw_rom(1326);
     when "010100101111" => data <= saw_rom(1327);
     when "010100110000" => data <= saw_rom(1328);
     when "010100110001" => data <= saw_rom(1329);
     when "010100110010" => data <= saw_rom(1330);
     when "010100110011" => data <= saw_rom(1331);
     when "010100110100" => data <= saw_rom(1332);
     when "010100110101" => data <= saw_rom(1333);
     when "010100110110" => data <= saw_rom(1334);
     when "010100110111" => data <= saw_rom(1335);
     when "010100111000" => data <= saw_rom(1336);
     when "010100111001" => data <= saw_rom(1337);
     when "010100111010" => data <= saw_rom(1338);
     when "010100111011" => data <= saw_rom(1339);
     when "010100111100" => data <= saw_rom(1340);
     when "010100111101" => data <= saw_rom(1341);
     when "010100111110" => data <= saw_rom(1342);
     when "010100111111" => data <= saw_rom(1343);
     when "010101000000" => data <= saw_rom(1344);
     when "010101000001" => data <= saw_rom(1345);
     when "010101000010" => data <= saw_rom(1346);
     when "010101000011" => data <= saw_rom(1347);
     when "010101000100" => data <= saw_rom(1348);
     when "010101000101" => data <= saw_rom(1349);
     when "010101000110" => data <= saw_rom(1350);
     when "010101000111" => data <= saw_rom(1351);
     when "010101001000" => data <= saw_rom(1352);
     when "010101001001" => data <= saw_rom(1353);
     when "010101001010" => data <= saw_rom(1354);
     when "010101001011" => data <= saw_rom(1355);
     when "010101001100" => data <= saw_rom(1356);
     when "010101001101" => data <= saw_rom(1357);
     when "010101001110" => data <= saw_rom(1358);
     when "010101001111" => data <= saw_rom(1359);
     when "010101010000" => data <= saw_rom(1360);
     when "010101010001" => data <= saw_rom(1361);
     when "010101010010" => data <= saw_rom(1362);
     when "010101010011" => data <= saw_rom(1363);
     when "010101010100" => data <= saw_rom(1364);
     when "010101010101" => data <= saw_rom(1365);
     when "010101010110" => data <= saw_rom(1366);
     when "010101010111" => data <= saw_rom(1367);
     when "010101011000" => data <= saw_rom(1368);
     when "010101011001" => data <= saw_rom(1369);
     when "010101011010" => data <= saw_rom(1370);
     when "010101011011" => data <= saw_rom(1371);
     when "010101011100" => data <= saw_rom(1372);
     when "010101011101" => data <= saw_rom(1373);
     when "010101011110" => data <= saw_rom(1374);
     when "010101011111" => data <= saw_rom(1375);
     when "010101100000" => data <= saw_rom(1376);
     when "010101100001" => data <= saw_rom(1377);
     when "010101100010" => data <= saw_rom(1378);
     when "010101100011" => data <= saw_rom(1379);
     when "010101100100" => data <= saw_rom(1380);
     when "010101100101" => data <= saw_rom(1381);
     when "010101100110" => data <= saw_rom(1382);
     when "010101100111" => data <= saw_rom(1383);
     when "010101101000" => data <= saw_rom(1384);
     when "010101101001" => data <= saw_rom(1385);
     when "010101101010" => data <= saw_rom(1386);
     when "010101101011" => data <= saw_rom(1387);
     when "010101101100" => data <= saw_rom(1388);
     when "010101101101" => data <= saw_rom(1389);
     when "010101101110" => data <= saw_rom(1390);
     when "010101101111" => data <= saw_rom(1391);
     when "010101110000" => data <= saw_rom(1392);
     when "010101110001" => data <= saw_rom(1393);
     when "010101110010" => data <= saw_rom(1394);
     when "010101110011" => data <= saw_rom(1395);
     when "010101110100" => data <= saw_rom(1396);
     when "010101110101" => data <= saw_rom(1397);
     when "010101110110" => data <= saw_rom(1398);
     when "010101110111" => data <= saw_rom(1399);
     when "010101111000" => data <= saw_rom(1400);
     when "010101111001" => data <= saw_rom(1401);
     when "010101111010" => data <= saw_rom(1402);
     when "010101111011" => data <= saw_rom(1403);
     when "010101111100" => data <= saw_rom(1404);
     when "010101111101" => data <= saw_rom(1405);
     when "010101111110" => data <= saw_rom(1406);
     when "010101111111" => data <= saw_rom(1407);
     when "010110000000" => data <= saw_rom(1408);
     when "010110000001" => data <= saw_rom(1409);
     when "010110000010" => data <= saw_rom(1410);
     when "010110000011" => data <= saw_rom(1411);
     when "010110000100" => data <= saw_rom(1412);
     when "010110000101" => data <= saw_rom(1413);
     when "010110000110" => data <= saw_rom(1414);
     when "010110000111" => data <= saw_rom(1415);
     when "010110001000" => data <= saw_rom(1416);
     when "010110001001" => data <= saw_rom(1417);
     when "010110001010" => data <= saw_rom(1418);
     when "010110001011" => data <= saw_rom(1419);
     when "010110001100" => data <= saw_rom(1420);
     when "010110001101" => data <= saw_rom(1421);
     when "010110001110" => data <= saw_rom(1422);
     when "010110001111" => data <= saw_rom(1423);
     when "010110010000" => data <= saw_rom(1424);
     when "010110010001" => data <= saw_rom(1425);
     when "010110010010" => data <= saw_rom(1426);
     when "010110010011" => data <= saw_rom(1427);
     when "010110010100" => data <= saw_rom(1428);
     when "010110010101" => data <= saw_rom(1429);
     when "010110010110" => data <= saw_rom(1430);
     when "010110010111" => data <= saw_rom(1431);
     when "010110011000" => data <= saw_rom(1432);
     when "010110011001" => data <= saw_rom(1433);
     when "010110011010" => data <= saw_rom(1434);
     when "010110011011" => data <= saw_rom(1435);
     when "010110011100" => data <= saw_rom(1436);
     when "010110011101" => data <= saw_rom(1437);
     when "010110011110" => data <= saw_rom(1438);
     when "010110011111" => data <= saw_rom(1439);
     when "010110100000" => data <= saw_rom(1440);
     when "010110100001" => data <= saw_rom(1441);
     when "010110100010" => data <= saw_rom(1442);
     when "010110100011" => data <= saw_rom(1443);
     when "010110100100" => data <= saw_rom(1444);
     when "010110100101" => data <= saw_rom(1445);
     when "010110100110" => data <= saw_rom(1446);
     when "010110100111" => data <= saw_rom(1447);
     when "010110101000" => data <= saw_rom(1448);
     when "010110101001" => data <= saw_rom(1449);
     when "010110101010" => data <= saw_rom(1450);
     when "010110101011" => data <= saw_rom(1451);
     when "010110101100" => data <= saw_rom(1452);
     when "010110101101" => data <= saw_rom(1453);
     when "010110101110" => data <= saw_rom(1454);
     when "010110101111" => data <= saw_rom(1455);
     when "010110110000" => data <= saw_rom(1456);
     when "010110110001" => data <= saw_rom(1457);
     when "010110110010" => data <= saw_rom(1458);
     when "010110110011" => data <= saw_rom(1459);
     when "010110110100" => data <= saw_rom(1460);
     when "010110110101" => data <= saw_rom(1461);
     when "010110110110" => data <= saw_rom(1462);
     when "010110110111" => data <= saw_rom(1463);
     when "010110111000" => data <= saw_rom(1464);
     when "010110111001" => data <= saw_rom(1465);
     when "010110111010" => data <= saw_rom(1466);
     when "010110111011" => data <= saw_rom(1467);
     when "010110111100" => data <= saw_rom(1468);
     when "010110111101" => data <= saw_rom(1469);
     when "010110111110" => data <= saw_rom(1470);
     when "010110111111" => data <= saw_rom(1471);
     when "010111000000" => data <= saw_rom(1472);
     when "010111000001" => data <= saw_rom(1473);
     when "010111000010" => data <= saw_rom(1474);
     when "010111000011" => data <= saw_rom(1475);
     when "010111000100" => data <= saw_rom(1476);
     when "010111000101" => data <= saw_rom(1477);
     when "010111000110" => data <= saw_rom(1478);
     when "010111000111" => data <= saw_rom(1479);
     when "010111001000" => data <= saw_rom(1480);
     when "010111001001" => data <= saw_rom(1481);
     when "010111001010" => data <= saw_rom(1482);
     when "010111001011" => data <= saw_rom(1483);
     when "010111001100" => data <= saw_rom(1484);
     when "010111001101" => data <= saw_rom(1485);
     when "010111001110" => data <= saw_rom(1486);
     when "010111001111" => data <= saw_rom(1487);
     when "010111010000" => data <= saw_rom(1488);
     when "010111010001" => data <= saw_rom(1489);
     when "010111010010" => data <= saw_rom(1490);
     when "010111010011" => data <= saw_rom(1491);
     when "010111010100" => data <= saw_rom(1492);
     when "010111010101" => data <= saw_rom(1493);
     when "010111010110" => data <= saw_rom(1494);
     when "010111010111" => data <= saw_rom(1495);
     when "010111011000" => data <= saw_rom(1496);
     when "010111011001" => data <= saw_rom(1497);
     when "010111011010" => data <= saw_rom(1498);
     when "010111011011" => data <= saw_rom(1499);
     when "010111011100" => data <= saw_rom(1500);
     when "010111011101" => data <= saw_rom(1501);
     when "010111011110" => data <= saw_rom(1502);
     when "010111011111" => data <= saw_rom(1503);
     when "010111100000" => data <= saw_rom(1504);
     when "010111100001" => data <= saw_rom(1505);
     when "010111100010" => data <= saw_rom(1506);
     when "010111100011" => data <= saw_rom(1507);
     when "010111100100" => data <= saw_rom(1508);
     when "010111100101" => data <= saw_rom(1509);
     when "010111100110" => data <= saw_rom(1510);
     when "010111100111" => data <= saw_rom(1511);
     when "010111101000" => data <= saw_rom(1512);
     when "010111101001" => data <= saw_rom(1513);
     when "010111101010" => data <= saw_rom(1514);
     when "010111101011" => data <= saw_rom(1515);
     when "010111101100" => data <= saw_rom(1516);
     when "010111101101" => data <= saw_rom(1517);
     when "010111101110" => data <= saw_rom(1518);
     when "010111101111" => data <= saw_rom(1519);
     when "010111110000" => data <= saw_rom(1520);
     when "010111110001" => data <= saw_rom(1521);
     when "010111110010" => data <= saw_rom(1522);
     when "010111110011" => data <= saw_rom(1523);
     when "010111110100" => data <= saw_rom(1524);
     when "010111110101" => data <= saw_rom(1525);
     when "010111110110" => data <= saw_rom(1526);
     when "010111110111" => data <= saw_rom(1527);
     when "010111111000" => data <= saw_rom(1528);
     when "010111111001" => data <= saw_rom(1529);
     when "010111111010" => data <= saw_rom(1530);
     when "010111111011" => data <= saw_rom(1531);
     when "010111111100" => data <= saw_rom(1532);
     when "010111111101" => data <= saw_rom(1533);
     when "010111111110" => data <= saw_rom(1534);
     when "010111111111" => data <= saw_rom(1535);
     when "011000000000" => data <= saw_rom(1536);
     when "011000000001" => data <= saw_rom(1537);
     when "011000000010" => data <= saw_rom(1538);
     when "011000000011" => data <= saw_rom(1539);
     when "011000000100" => data <= saw_rom(1540);
     when "011000000101" => data <= saw_rom(1541);
     when "011000000110" => data <= saw_rom(1542);
     when "011000000111" => data <= saw_rom(1543);
     when "011000001000" => data <= saw_rom(1544);
     when "011000001001" => data <= saw_rom(1545);
     when "011000001010" => data <= saw_rom(1546);
     when "011000001011" => data <= saw_rom(1547);
     when "011000001100" => data <= saw_rom(1548);
     when "011000001101" => data <= saw_rom(1549);
     when "011000001110" => data <= saw_rom(1550);
     when "011000001111" => data <= saw_rom(1551);
     when "011000010000" => data <= saw_rom(1552);
     when "011000010001" => data <= saw_rom(1553);
     when "011000010010" => data <= saw_rom(1554);
     when "011000010011" => data <= saw_rom(1555);
     when "011000010100" => data <= saw_rom(1556);
     when "011000010101" => data <= saw_rom(1557);
     when "011000010110" => data <= saw_rom(1558);
     when "011000010111" => data <= saw_rom(1559);
     when "011000011000" => data <= saw_rom(1560);
     when "011000011001" => data <= saw_rom(1561);
     when "011000011010" => data <= saw_rom(1562);
     when "011000011011" => data <= saw_rom(1563);
     when "011000011100" => data <= saw_rom(1564);
     when "011000011101" => data <= saw_rom(1565);
     when "011000011110" => data <= saw_rom(1566);
     when "011000011111" => data <= saw_rom(1567);
     when "011000100000" => data <= saw_rom(1568);
     when "011000100001" => data <= saw_rom(1569);
     when "011000100010" => data <= saw_rom(1570);
     when "011000100011" => data <= saw_rom(1571);
     when "011000100100" => data <= saw_rom(1572);
     when "011000100101" => data <= saw_rom(1573);
     when "011000100110" => data <= saw_rom(1574);
     when "011000100111" => data <= saw_rom(1575);
     when "011000101000" => data <= saw_rom(1576);
     when "011000101001" => data <= saw_rom(1577);
     when "011000101010" => data <= saw_rom(1578);
     when "011000101011" => data <= saw_rom(1579);
     when "011000101100" => data <= saw_rom(1580);
     when "011000101101" => data <= saw_rom(1581);
     when "011000101110" => data <= saw_rom(1582);
     when "011000101111" => data <= saw_rom(1583);
     when "011000110000" => data <= saw_rom(1584);
     when "011000110001" => data <= saw_rom(1585);
     when "011000110010" => data <= saw_rom(1586);
     when "011000110011" => data <= saw_rom(1587);
     when "011000110100" => data <= saw_rom(1588);
     when "011000110101" => data <= saw_rom(1589);
     when "011000110110" => data <= saw_rom(1590);
     when "011000110111" => data <= saw_rom(1591);
     when "011000111000" => data <= saw_rom(1592);
     when "011000111001" => data <= saw_rom(1593);
     when "011000111010" => data <= saw_rom(1594);
     when "011000111011" => data <= saw_rom(1595);
     when "011000111100" => data <= saw_rom(1596);
     when "011000111101" => data <= saw_rom(1597);
     when "011000111110" => data <= saw_rom(1598);
     when "011000111111" => data <= saw_rom(1599);
     when "011001000000" => data <= saw_rom(1600);
     when "011001000001" => data <= saw_rom(1601);
     when "011001000010" => data <= saw_rom(1602);
     when "011001000011" => data <= saw_rom(1603);
     when "011001000100" => data <= saw_rom(1604);
     when "011001000101" => data <= saw_rom(1605);
     when "011001000110" => data <= saw_rom(1606);
     when "011001000111" => data <= saw_rom(1607);
     when "011001001000" => data <= saw_rom(1608);
     when "011001001001" => data <= saw_rom(1609);
     when "011001001010" => data <= saw_rom(1610);
     when "011001001011" => data <= saw_rom(1611);
     when "011001001100" => data <= saw_rom(1612);
     when "011001001101" => data <= saw_rom(1613);
     when "011001001110" => data <= saw_rom(1614);
     when "011001001111" => data <= saw_rom(1615);
     when "011001010000" => data <= saw_rom(1616);
     when "011001010001" => data <= saw_rom(1617);
     when "011001010010" => data <= saw_rom(1618);
     when "011001010011" => data <= saw_rom(1619);
     when "011001010100" => data <= saw_rom(1620);
     when "011001010101" => data <= saw_rom(1621);
     when "011001010110" => data <= saw_rom(1622);
     when "011001010111" => data <= saw_rom(1623);
     when "011001011000" => data <= saw_rom(1624);
     when "011001011001" => data <= saw_rom(1625);
     when "011001011010" => data <= saw_rom(1626);
     when "011001011011" => data <= saw_rom(1627);
     when "011001011100" => data <= saw_rom(1628);
     when "011001011101" => data <= saw_rom(1629);
     when "011001011110" => data <= saw_rom(1630);
     when "011001011111" => data <= saw_rom(1631);
     when "011001100000" => data <= saw_rom(1632);
     when "011001100001" => data <= saw_rom(1633);
     when "011001100010" => data <= saw_rom(1634);
     when "011001100011" => data <= saw_rom(1635);
     when "011001100100" => data <= saw_rom(1636);
     when "011001100101" => data <= saw_rom(1637);
     when "011001100110" => data <= saw_rom(1638);
     when "011001100111" => data <= saw_rom(1639);
     when "011001101000" => data <= saw_rom(1640);
     when "011001101001" => data <= saw_rom(1641);
     when "011001101010" => data <= saw_rom(1642);
     when "011001101011" => data <= saw_rom(1643);
     when "011001101100" => data <= saw_rom(1644);
     when "011001101101" => data <= saw_rom(1645);
     when "011001101110" => data <= saw_rom(1646);
     when "011001101111" => data <= saw_rom(1647);
     when "011001110000" => data <= saw_rom(1648);
     when "011001110001" => data <= saw_rom(1649);
     when "011001110010" => data <= saw_rom(1650);
     when "011001110011" => data <= saw_rom(1651);
     when "011001110100" => data <= saw_rom(1652);
     when "011001110101" => data <= saw_rom(1653);
     when "011001110110" => data <= saw_rom(1654);
     when "011001110111" => data <= saw_rom(1655);
     when "011001111000" => data <= saw_rom(1656);
     when "011001111001" => data <= saw_rom(1657);
     when "011001111010" => data <= saw_rom(1658);
     when "011001111011" => data <= saw_rom(1659);
     when "011001111100" => data <= saw_rom(1660);
     when "011001111101" => data <= saw_rom(1661);
     when "011001111110" => data <= saw_rom(1662);
     when "011001111111" => data <= saw_rom(1663);
     when "011010000000" => data <= saw_rom(1664);
     when "011010000001" => data <= saw_rom(1665);
     when "011010000010" => data <= saw_rom(1666);
     when "011010000011" => data <= saw_rom(1667);
     when "011010000100" => data <= saw_rom(1668);
     when "011010000101" => data <= saw_rom(1669);
     when "011010000110" => data <= saw_rom(1670);
     when "011010000111" => data <= saw_rom(1671);
     when "011010001000" => data <= saw_rom(1672);
     when "011010001001" => data <= saw_rom(1673);
     when "011010001010" => data <= saw_rom(1674);
     when "011010001011" => data <= saw_rom(1675);
     when "011010001100" => data <= saw_rom(1676);
     when "011010001101" => data <= saw_rom(1677);
     when "011010001110" => data <= saw_rom(1678);
     when "011010001111" => data <= saw_rom(1679);
     when "011010010000" => data <= saw_rom(1680);
     when "011010010001" => data <= saw_rom(1681);
     when "011010010010" => data <= saw_rom(1682);
     when "011010010011" => data <= saw_rom(1683);
     when "011010010100" => data <= saw_rom(1684);
     when "011010010101" => data <= saw_rom(1685);
     when "011010010110" => data <= saw_rom(1686);
     when "011010010111" => data <= saw_rom(1687);
     when "011010011000" => data <= saw_rom(1688);
     when "011010011001" => data <= saw_rom(1689);
     when "011010011010" => data <= saw_rom(1690);
     when "011010011011" => data <= saw_rom(1691);
     when "011010011100" => data <= saw_rom(1692);
     when "011010011101" => data <= saw_rom(1693);
     when "011010011110" => data <= saw_rom(1694);
     when "011010011111" => data <= saw_rom(1695);
     when "011010100000" => data <= saw_rom(1696);
     when "011010100001" => data <= saw_rom(1697);
     when "011010100010" => data <= saw_rom(1698);
     when "011010100011" => data <= saw_rom(1699);
     when "011010100100" => data <= saw_rom(1700);
     when "011010100101" => data <= saw_rom(1701);
     when "011010100110" => data <= saw_rom(1702);
     when "011010100111" => data <= saw_rom(1703);
     when "011010101000" => data <= saw_rom(1704);
     when "011010101001" => data <= saw_rom(1705);
     when "011010101010" => data <= saw_rom(1706);
     when "011010101011" => data <= saw_rom(1707);
     when "011010101100" => data <= saw_rom(1708);
     when "011010101101" => data <= saw_rom(1709);
     when "011010101110" => data <= saw_rom(1710);
     when "011010101111" => data <= saw_rom(1711);
     when "011010110000" => data <= saw_rom(1712);
     when "011010110001" => data <= saw_rom(1713);
     when "011010110010" => data <= saw_rom(1714);
     when "011010110011" => data <= saw_rom(1715);
     when "011010110100" => data <= saw_rom(1716);
     when "011010110101" => data <= saw_rom(1717);
     when "011010110110" => data <= saw_rom(1718);
     when "011010110111" => data <= saw_rom(1719);
     when "011010111000" => data <= saw_rom(1720);
     when "011010111001" => data <= saw_rom(1721);
     when "011010111010" => data <= saw_rom(1722);
     when "011010111011" => data <= saw_rom(1723);
     when "011010111100" => data <= saw_rom(1724);
     when "011010111101" => data <= saw_rom(1725);
     when "011010111110" => data <= saw_rom(1726);
     when "011010111111" => data <= saw_rom(1727);
     when "011011000000" => data <= saw_rom(1728);
     when "011011000001" => data <= saw_rom(1729);
     when "011011000010" => data <= saw_rom(1730);
     when "011011000011" => data <= saw_rom(1731);
     when "011011000100" => data <= saw_rom(1732);
     when "011011000101" => data <= saw_rom(1733);
     when "011011000110" => data <= saw_rom(1734);
     when "011011000111" => data <= saw_rom(1735);
     when "011011001000" => data <= saw_rom(1736);
     when "011011001001" => data <= saw_rom(1737);
     when "011011001010" => data <= saw_rom(1738);
     when "011011001011" => data <= saw_rom(1739);
     when "011011001100" => data <= saw_rom(1740);
     when "011011001101" => data <= saw_rom(1741);
     when "011011001110" => data <= saw_rom(1742);
     when "011011001111" => data <= saw_rom(1743);
     when "011011010000" => data <= saw_rom(1744);
     when "011011010001" => data <= saw_rom(1745);
     when "011011010010" => data <= saw_rom(1746);
     when "011011010011" => data <= saw_rom(1747);
     when "011011010100" => data <= saw_rom(1748);
     when "011011010101" => data <= saw_rom(1749);
     when "011011010110" => data <= saw_rom(1750);
     when "011011010111" => data <= saw_rom(1751);
     when "011011011000" => data <= saw_rom(1752);
     when "011011011001" => data <= saw_rom(1753);
     when "011011011010" => data <= saw_rom(1754);
     when "011011011011" => data <= saw_rom(1755);
     when "011011011100" => data <= saw_rom(1756);
     when "011011011101" => data <= saw_rom(1757);
     when "011011011110" => data <= saw_rom(1758);
     when "011011011111" => data <= saw_rom(1759);
     when "011011100000" => data <= saw_rom(1760);
     when "011011100001" => data <= saw_rom(1761);
     when "011011100010" => data <= saw_rom(1762);
     when "011011100011" => data <= saw_rom(1763);
     when "011011100100" => data <= saw_rom(1764);
     when "011011100101" => data <= saw_rom(1765);
     when "011011100110" => data <= saw_rom(1766);
     when "011011100111" => data <= saw_rom(1767);
     when "011011101000" => data <= saw_rom(1768);
     when "011011101001" => data <= saw_rom(1769);
     when "011011101010" => data <= saw_rom(1770);
     when "011011101011" => data <= saw_rom(1771);
     when "011011101100" => data <= saw_rom(1772);
     when "011011101101" => data <= saw_rom(1773);
     when "011011101110" => data <= saw_rom(1774);
     when "011011101111" => data <= saw_rom(1775);
     when "011011110000" => data <= saw_rom(1776);
     when "011011110001" => data <= saw_rom(1777);
     when "011011110010" => data <= saw_rom(1778);
     when "011011110011" => data <= saw_rom(1779);
     when "011011110100" => data <= saw_rom(1780);
     when "011011110101" => data <= saw_rom(1781);
     when "011011110110" => data <= saw_rom(1782);
     when "011011110111" => data <= saw_rom(1783);
     when "011011111000" => data <= saw_rom(1784);
     when "011011111001" => data <= saw_rom(1785);
     when "011011111010" => data <= saw_rom(1786);
     when "011011111011" => data <= saw_rom(1787);
     when "011011111100" => data <= saw_rom(1788);
     when "011011111101" => data <= saw_rom(1789);
     when "011011111110" => data <= saw_rom(1790);
     when "011011111111" => data <= saw_rom(1791);
     when "011100000000" => data <= saw_rom(1792);
     when "011100000001" => data <= saw_rom(1793);
     when "011100000010" => data <= saw_rom(1794);
     when "011100000011" => data <= saw_rom(1795);
     when "011100000100" => data <= saw_rom(1796);
     when "011100000101" => data <= saw_rom(1797);
     when "011100000110" => data <= saw_rom(1798);
     when "011100000111" => data <= saw_rom(1799);
     when "011100001000" => data <= saw_rom(1800);
     when "011100001001" => data <= saw_rom(1801);
     when "011100001010" => data <= saw_rom(1802);
     when "011100001011" => data <= saw_rom(1803);
     when "011100001100" => data <= saw_rom(1804);
     when "011100001101" => data <= saw_rom(1805);
     when "011100001110" => data <= saw_rom(1806);
     when "011100001111" => data <= saw_rom(1807);
     when "011100010000" => data <= saw_rom(1808);
     when "011100010001" => data <= saw_rom(1809);
     when "011100010010" => data <= saw_rom(1810);
     when "011100010011" => data <= saw_rom(1811);
     when "011100010100" => data <= saw_rom(1812);
     when "011100010101" => data <= saw_rom(1813);
     when "011100010110" => data <= saw_rom(1814);
     when "011100010111" => data <= saw_rom(1815);
     when "011100011000" => data <= saw_rom(1816);
     when "011100011001" => data <= saw_rom(1817);
     when "011100011010" => data <= saw_rom(1818);
     when "011100011011" => data <= saw_rom(1819);
     when "011100011100" => data <= saw_rom(1820);
     when "011100011101" => data <= saw_rom(1821);
     when "011100011110" => data <= saw_rom(1822);
     when "011100011111" => data <= saw_rom(1823);
     when "011100100000" => data <= saw_rom(1824);
     when "011100100001" => data <= saw_rom(1825);
     when "011100100010" => data <= saw_rom(1826);
     when "011100100011" => data <= saw_rom(1827);
     when "011100100100" => data <= saw_rom(1828);
     when "011100100101" => data <= saw_rom(1829);
     when "011100100110" => data <= saw_rom(1830);
     when "011100100111" => data <= saw_rom(1831);
     when "011100101000" => data <= saw_rom(1832);
     when "011100101001" => data <= saw_rom(1833);
     when "011100101010" => data <= saw_rom(1834);
     when "011100101011" => data <= saw_rom(1835);
     when "011100101100" => data <= saw_rom(1836);
     when "011100101101" => data <= saw_rom(1837);
     when "011100101110" => data <= saw_rom(1838);
     when "011100101111" => data <= saw_rom(1839);
     when "011100110000" => data <= saw_rom(1840);
     when "011100110001" => data <= saw_rom(1841);
     when "011100110010" => data <= saw_rom(1842);
     when "011100110011" => data <= saw_rom(1843);
     when "011100110100" => data <= saw_rom(1844);
     when "011100110101" => data <= saw_rom(1845);
     when "011100110110" => data <= saw_rom(1846);
     when "011100110111" => data <= saw_rom(1847);
     when "011100111000" => data <= saw_rom(1848);
     when "011100111001" => data <= saw_rom(1849);
     when "011100111010" => data <= saw_rom(1850);
     when "011100111011" => data <= saw_rom(1851);
     when "011100111100" => data <= saw_rom(1852);
     when "011100111101" => data <= saw_rom(1853);
     when "011100111110" => data <= saw_rom(1854);
     when "011100111111" => data <= saw_rom(1855);
     when "011101000000" => data <= saw_rom(1856);
     when "011101000001" => data <= saw_rom(1857);
     when "011101000010" => data <= saw_rom(1858);
     when "011101000011" => data <= saw_rom(1859);
     when "011101000100" => data <= saw_rom(1860);
     when "011101000101" => data <= saw_rom(1861);
     when "011101000110" => data <= saw_rom(1862);
     when "011101000111" => data <= saw_rom(1863);
     when "011101001000" => data <= saw_rom(1864);
     when "011101001001" => data <= saw_rom(1865);
     when "011101001010" => data <= saw_rom(1866);
     when "011101001011" => data <= saw_rom(1867);
     when "011101001100" => data <= saw_rom(1868);
     when "011101001101" => data <= saw_rom(1869);
     when "011101001110" => data <= saw_rom(1870);
     when "011101001111" => data <= saw_rom(1871);
     when "011101010000" => data <= saw_rom(1872);
     when "011101010001" => data <= saw_rom(1873);
     when "011101010010" => data <= saw_rom(1874);
     when "011101010011" => data <= saw_rom(1875);
     when "011101010100" => data <= saw_rom(1876);
     when "011101010101" => data <= saw_rom(1877);
     when "011101010110" => data <= saw_rom(1878);
     when "011101010111" => data <= saw_rom(1879);
     when "011101011000" => data <= saw_rom(1880);
     when "011101011001" => data <= saw_rom(1881);
     when "011101011010" => data <= saw_rom(1882);
     when "011101011011" => data <= saw_rom(1883);
     when "011101011100" => data <= saw_rom(1884);
     when "011101011101" => data <= saw_rom(1885);
     when "011101011110" => data <= saw_rom(1886);
     when "011101011111" => data <= saw_rom(1887);
     when "011101100000" => data <= saw_rom(1888);
     when "011101100001" => data <= saw_rom(1889);
     when "011101100010" => data <= saw_rom(1890);
     when "011101100011" => data <= saw_rom(1891);
     when "011101100100" => data <= saw_rom(1892);
     when "011101100101" => data <= saw_rom(1893);
     when "011101100110" => data <= saw_rom(1894);
     when "011101100111" => data <= saw_rom(1895);
     when "011101101000" => data <= saw_rom(1896);
     when "011101101001" => data <= saw_rom(1897);
     when "011101101010" => data <= saw_rom(1898);
     when "011101101011" => data <= saw_rom(1899);
     when "011101101100" => data <= saw_rom(1900);
     when "011101101101" => data <= saw_rom(1901);
     when "011101101110" => data <= saw_rom(1902);
     when "011101101111" => data <= saw_rom(1903);
     when "011101110000" => data <= saw_rom(1904);
     when "011101110001" => data <= saw_rom(1905);
     when "011101110010" => data <= saw_rom(1906);
     when "011101110011" => data <= saw_rom(1907);
     when "011101110100" => data <= saw_rom(1908);
     when "011101110101" => data <= saw_rom(1909);
     when "011101110110" => data <= saw_rom(1910);
     when "011101110111" => data <= saw_rom(1911);
     when "011101111000" => data <= saw_rom(1912);
     when "011101111001" => data <= saw_rom(1913);
     when "011101111010" => data <= saw_rom(1914);
     when "011101111011" => data <= saw_rom(1915);
     when "011101111100" => data <= saw_rom(1916);
     when "011101111101" => data <= saw_rom(1917);
     when "011101111110" => data <= saw_rom(1918);
     when "011101111111" => data <= saw_rom(1919);
     when "011110000000" => data <= saw_rom(1920);
     when "011110000001" => data <= saw_rom(1921);
     when "011110000010" => data <= saw_rom(1922);
     when "011110000011" => data <= saw_rom(1923);
     when "011110000100" => data <= saw_rom(1924);
     when "011110000101" => data <= saw_rom(1925);
     when "011110000110" => data <= saw_rom(1926);
     when "011110000111" => data <= saw_rom(1927);
     when "011110001000" => data <= saw_rom(1928);
     when "011110001001" => data <= saw_rom(1929);
     when "011110001010" => data <= saw_rom(1930);
     when "011110001011" => data <= saw_rom(1931);
     when "011110001100" => data <= saw_rom(1932);
     when "011110001101" => data <= saw_rom(1933);
     when "011110001110" => data <= saw_rom(1934);
     when "011110001111" => data <= saw_rom(1935);
     when "011110010000" => data <= saw_rom(1936);
     when "011110010001" => data <= saw_rom(1937);
     when "011110010010" => data <= saw_rom(1938);
     when "011110010011" => data <= saw_rom(1939);
     when "011110010100" => data <= saw_rom(1940);
     when "011110010101" => data <= saw_rom(1941);
     when "011110010110" => data <= saw_rom(1942);
     when "011110010111" => data <= saw_rom(1943);
     when "011110011000" => data <= saw_rom(1944);
     when "011110011001" => data <= saw_rom(1945);
     when "011110011010" => data <= saw_rom(1946);
     when "011110011011" => data <= saw_rom(1947);
     when "011110011100" => data <= saw_rom(1948);
     when "011110011101" => data <= saw_rom(1949);
     when "011110011110" => data <= saw_rom(1950);
     when "011110011111" => data <= saw_rom(1951);
     when "011110100000" => data <= saw_rom(1952);
     when "011110100001" => data <= saw_rom(1953);
     when "011110100010" => data <= saw_rom(1954);
     when "011110100011" => data <= saw_rom(1955);
     when "011110100100" => data <= saw_rom(1956);
     when "011110100101" => data <= saw_rom(1957);
     when "011110100110" => data <= saw_rom(1958);
     when "011110100111" => data <= saw_rom(1959);
     when "011110101000" => data <= saw_rom(1960);
     when "011110101001" => data <= saw_rom(1961);
     when "011110101010" => data <= saw_rom(1962);
     when "011110101011" => data <= saw_rom(1963);
     when "011110101100" => data <= saw_rom(1964);
     when "011110101101" => data <= saw_rom(1965);
     when "011110101110" => data <= saw_rom(1966);
     when "011110101111" => data <= saw_rom(1967);
     when "011110110000" => data <= saw_rom(1968);
     when "011110110001" => data <= saw_rom(1969);
     when "011110110010" => data <= saw_rom(1970);
     when "011110110011" => data <= saw_rom(1971);
     when "011110110100" => data <= saw_rom(1972);
     when "011110110101" => data <= saw_rom(1973);
     when "011110110110" => data <= saw_rom(1974);
     when "011110110111" => data <= saw_rom(1975);
     when "011110111000" => data <= saw_rom(1976);
     when "011110111001" => data <= saw_rom(1977);
     when "011110111010" => data <= saw_rom(1978);
     when "011110111011" => data <= saw_rom(1979);
     when "011110111100" => data <= saw_rom(1980);
     when "011110111101" => data <= saw_rom(1981);
     when "011110111110" => data <= saw_rom(1982);
     when "011110111111" => data <= saw_rom(1983);
     when "011111000000" => data <= saw_rom(1984);
     when "011111000001" => data <= saw_rom(1985);
     when "011111000010" => data <= saw_rom(1986);
     when "011111000011" => data <= saw_rom(1987);
     when "011111000100" => data <= saw_rom(1988);
     when "011111000101" => data <= saw_rom(1989);
     when "011111000110" => data <= saw_rom(1990);
     when "011111000111" => data <= saw_rom(1991);
     when "011111001000" => data <= saw_rom(1992);
     when "011111001001" => data <= saw_rom(1993);
     when "011111001010" => data <= saw_rom(1994);
     when "011111001011" => data <= saw_rom(1995);
     when "011111001100" => data <= saw_rom(1996);
     when "011111001101" => data <= saw_rom(1997);
     when "011111001110" => data <= saw_rom(1998);
     when "011111001111" => data <= saw_rom(1999);
     when "011111010000" => data <= saw_rom(2000);
     when "011111010001" => data <= saw_rom(2001);
     when "011111010010" => data <= saw_rom(2002);
     when "011111010011" => data <= saw_rom(2003);
     when "011111010100" => data <= saw_rom(2004);
     when "011111010101" => data <= saw_rom(2005);
     when "011111010110" => data <= saw_rom(2006);
     when "011111010111" => data <= saw_rom(2007);
     when "011111011000" => data <= saw_rom(2008);
     when "011111011001" => data <= saw_rom(2009);
     when "011111011010" => data <= saw_rom(2010);
     when "011111011011" => data <= saw_rom(2011);
     when "011111011100" => data <= saw_rom(2012);
     when "011111011101" => data <= saw_rom(2013);
     when "011111011110" => data <= saw_rom(2014);
     when "011111011111" => data <= saw_rom(2015);
     when "011111100000" => data <= saw_rom(2016);
     when "011111100001" => data <= saw_rom(2017);
     when "011111100010" => data <= saw_rom(2018);
     when "011111100011" => data <= saw_rom(2019);
     when "011111100100" => data <= saw_rom(2020);
     when "011111100101" => data <= saw_rom(2021);
     when "011111100110" => data <= saw_rom(2022);
     when "011111100111" => data <= saw_rom(2023);
     when "011111101000" => data <= saw_rom(2024);
     when "011111101001" => data <= saw_rom(2025);
     when "011111101010" => data <= saw_rom(2026);
     when "011111101011" => data <= saw_rom(2027);
     when "011111101100" => data <= saw_rom(2028);
     when "011111101101" => data <= saw_rom(2029);
     when "011111101110" => data <= saw_rom(2030);
     when "011111101111" => data <= saw_rom(2031);
     when "011111110000" => data <= saw_rom(2032);
     when "011111110001" => data <= saw_rom(2033);
     when "011111110010" => data <= saw_rom(2034);
     when "011111110011" => data <= saw_rom(2035);
     when "011111110100" => data <= saw_rom(2036);
     when "011111110101" => data <= saw_rom(2037);
     when "011111110110" => data <= saw_rom(2038);
     when "011111110111" => data <= saw_rom(2039);
     when "011111111000" => data <= saw_rom(2040);
     when "011111111001" => data <= saw_rom(2041);
     when "011111111010" => data <= saw_rom(2042);
     when "011111111011" => data <= saw_rom(2043);
     when "011111111100" => data <= saw_rom(2044);
     when "011111111101" => data <= saw_rom(2045);
     when "011111111110" => data <= saw_rom(2046);
     when "011111111111" => data <= saw_rom(2047);
     when "100000000000" => data <= saw_rom(2048);
     when "100000000001" => data <= saw_rom(2049);
     when "100000000010" => data <= saw_rom(2050);
     when "100000000011" => data <= saw_rom(2051);
     when "100000000100" => data <= saw_rom(2052);
     when "100000000101" => data <= saw_rom(2053);
     when "100000000110" => data <= saw_rom(2054);
     when "100000000111" => data <= saw_rom(2055);
     when "100000001000" => data <= saw_rom(2056);
     when "100000001001" => data <= saw_rom(2057);
     when "100000001010" => data <= saw_rom(2058);
     when "100000001011" => data <= saw_rom(2059);
     when "100000001100" => data <= saw_rom(2060);
     when "100000001101" => data <= saw_rom(2061);
     when "100000001110" => data <= saw_rom(2062);
     when "100000001111" => data <= saw_rom(2063);
     when "100000010000" => data <= saw_rom(2064);
     when "100000010001" => data <= saw_rom(2065);
     when "100000010010" => data <= saw_rom(2066);
     when "100000010011" => data <= saw_rom(2067);
     when "100000010100" => data <= saw_rom(2068);
     when "100000010101" => data <= saw_rom(2069);
     when "100000010110" => data <= saw_rom(2070);
     when "100000010111" => data <= saw_rom(2071);
     when "100000011000" => data <= saw_rom(2072);
     when "100000011001" => data <= saw_rom(2073);
     when "100000011010" => data <= saw_rom(2074);
     when "100000011011" => data <= saw_rom(2075);
     when "100000011100" => data <= saw_rom(2076);
     when "100000011101" => data <= saw_rom(2077);
     when "100000011110" => data <= saw_rom(2078);
     when "100000011111" => data <= saw_rom(2079);
     when "100000100000" => data <= saw_rom(2080);
     when "100000100001" => data <= saw_rom(2081);
     when "100000100010" => data <= saw_rom(2082);
     when "100000100011" => data <= saw_rom(2083);
     when "100000100100" => data <= saw_rom(2084);
     when "100000100101" => data <= saw_rom(2085);
     when "100000100110" => data <= saw_rom(2086);
     when "100000100111" => data <= saw_rom(2087);
     when "100000101000" => data <= saw_rom(2088);
     when "100000101001" => data <= saw_rom(2089);
     when "100000101010" => data <= saw_rom(2090);
     when "100000101011" => data <= saw_rom(2091);
     when "100000101100" => data <= saw_rom(2092);
     when "100000101101" => data <= saw_rom(2093);
     when "100000101110" => data <= saw_rom(2094);
     when "100000101111" => data <= saw_rom(2095);
     when "100000110000" => data <= saw_rom(2096);
     when "100000110001" => data <= saw_rom(2097);
     when "100000110010" => data <= saw_rom(2098);
     when "100000110011" => data <= saw_rom(2099);
     when "100000110100" => data <= saw_rom(2100);
     when "100000110101" => data <= saw_rom(2101);
     when "100000110110" => data <= saw_rom(2102);
     when "100000110111" => data <= saw_rom(2103);
     when "100000111000" => data <= saw_rom(2104);
     when "100000111001" => data <= saw_rom(2105);
     when "100000111010" => data <= saw_rom(2106);
     when "100000111011" => data <= saw_rom(2107);
     when "100000111100" => data <= saw_rom(2108);
     when "100000111101" => data <= saw_rom(2109);
     when "100000111110" => data <= saw_rom(2110);
     when "100000111111" => data <= saw_rom(2111);
     when "100001000000" => data <= saw_rom(2112);
     when "100001000001" => data <= saw_rom(2113);
     when "100001000010" => data <= saw_rom(2114);
     when "100001000011" => data <= saw_rom(2115);
     when "100001000100" => data <= saw_rom(2116);
     when "100001000101" => data <= saw_rom(2117);
     when "100001000110" => data <= saw_rom(2118);
     when "100001000111" => data <= saw_rom(2119);
     when "100001001000" => data <= saw_rom(2120);
     when "100001001001" => data <= saw_rom(2121);
     when "100001001010" => data <= saw_rom(2122);
     when "100001001011" => data <= saw_rom(2123);
     when "100001001100" => data <= saw_rom(2124);
     when "100001001101" => data <= saw_rom(2125);
     when "100001001110" => data <= saw_rom(2126);
     when "100001001111" => data <= saw_rom(2127);
     when "100001010000" => data <= saw_rom(2128);
     when "100001010001" => data <= saw_rom(2129);
     when "100001010010" => data <= saw_rom(2130);
     when "100001010011" => data <= saw_rom(2131);
     when "100001010100" => data <= saw_rom(2132);
     when "100001010101" => data <= saw_rom(2133);
     when "100001010110" => data <= saw_rom(2134);
     when "100001010111" => data <= saw_rom(2135);
     when "100001011000" => data <= saw_rom(2136);
     when "100001011001" => data <= saw_rom(2137);
     when "100001011010" => data <= saw_rom(2138);
     when "100001011011" => data <= saw_rom(2139);
     when "100001011100" => data <= saw_rom(2140);
     when "100001011101" => data <= saw_rom(2141);
     when "100001011110" => data <= saw_rom(2142);
     when "100001011111" => data <= saw_rom(2143);
     when "100001100000" => data <= saw_rom(2144);
     when "100001100001" => data <= saw_rom(2145);
     when "100001100010" => data <= saw_rom(2146);
     when "100001100011" => data <= saw_rom(2147);
     when "100001100100" => data <= saw_rom(2148);
     when "100001100101" => data <= saw_rom(2149);
     when "100001100110" => data <= saw_rom(2150);
     when "100001100111" => data <= saw_rom(2151);
     when "100001101000" => data <= saw_rom(2152);
     when "100001101001" => data <= saw_rom(2153);
     when "100001101010" => data <= saw_rom(2154);
     when "100001101011" => data <= saw_rom(2155);
     when "100001101100" => data <= saw_rom(2156);
     when "100001101101" => data <= saw_rom(2157);
     when "100001101110" => data <= saw_rom(2158);
     when "100001101111" => data <= saw_rom(2159);
     when "100001110000" => data <= saw_rom(2160);
     when "100001110001" => data <= saw_rom(2161);
     when "100001110010" => data <= saw_rom(2162);
     when "100001110011" => data <= saw_rom(2163);
     when "100001110100" => data <= saw_rom(2164);
     when "100001110101" => data <= saw_rom(2165);
     when "100001110110" => data <= saw_rom(2166);
     when "100001110111" => data <= saw_rom(2167);
     when "100001111000" => data <= saw_rom(2168);
     when "100001111001" => data <= saw_rom(2169);
     when "100001111010" => data <= saw_rom(2170);
     when "100001111011" => data <= saw_rom(2171);
     when "100001111100" => data <= saw_rom(2172);
     when "100001111101" => data <= saw_rom(2173);
     when "100001111110" => data <= saw_rom(2174);
     when "100001111111" => data <= saw_rom(2175);
     when "100010000000" => data <= saw_rom(2176);
     when "100010000001" => data <= saw_rom(2177);
     when "100010000010" => data <= saw_rom(2178);
     when "100010000011" => data <= saw_rom(2179);
     when "100010000100" => data <= saw_rom(2180);
     when "100010000101" => data <= saw_rom(2181);
     when "100010000110" => data <= saw_rom(2182);
     when "100010000111" => data <= saw_rom(2183);
     when "100010001000" => data <= saw_rom(2184);
     when "100010001001" => data <= saw_rom(2185);
     when "100010001010" => data <= saw_rom(2186);
     when "100010001011" => data <= saw_rom(2187);
     when "100010001100" => data <= saw_rom(2188);
     when "100010001101" => data <= saw_rom(2189);
     when "100010001110" => data <= saw_rom(2190);
     when "100010001111" => data <= saw_rom(2191);
     when "100010010000" => data <= saw_rom(2192);
     when "100010010001" => data <= saw_rom(2193);
     when "100010010010" => data <= saw_rom(2194);
     when "100010010011" => data <= saw_rom(2195);
     when "100010010100" => data <= saw_rom(2196);
     when "100010010101" => data <= saw_rom(2197);
     when "100010010110" => data <= saw_rom(2198);
     when "100010010111" => data <= saw_rom(2199);
     when "100010011000" => data <= saw_rom(2200);
     when "100010011001" => data <= saw_rom(2201);
     when "100010011010" => data <= saw_rom(2202);
     when "100010011011" => data <= saw_rom(2203);
     when "100010011100" => data <= saw_rom(2204);
     when "100010011101" => data <= saw_rom(2205);
     when "100010011110" => data <= saw_rom(2206);
     when "100010011111" => data <= saw_rom(2207);
     when "100010100000" => data <= saw_rom(2208);
     when "100010100001" => data <= saw_rom(2209);
     when "100010100010" => data <= saw_rom(2210);
     when "100010100011" => data <= saw_rom(2211);
     when "100010100100" => data <= saw_rom(2212);
     when "100010100101" => data <= saw_rom(2213);
     when "100010100110" => data <= saw_rom(2214);
     when "100010100111" => data <= saw_rom(2215);
     when "100010101000" => data <= saw_rom(2216);
     when "100010101001" => data <= saw_rom(2217);
     when "100010101010" => data <= saw_rom(2218);
     when "100010101011" => data <= saw_rom(2219);
     when "100010101100" => data <= saw_rom(2220);
     when "100010101101" => data <= saw_rom(2221);
     when "100010101110" => data <= saw_rom(2222);
     when "100010101111" => data <= saw_rom(2223);
     when "100010110000" => data <= saw_rom(2224);
     when "100010110001" => data <= saw_rom(2225);
     when "100010110010" => data <= saw_rom(2226);
     when "100010110011" => data <= saw_rom(2227);
     when "100010110100" => data <= saw_rom(2228);
     when "100010110101" => data <= saw_rom(2229);
     when "100010110110" => data <= saw_rom(2230);
     when "100010110111" => data <= saw_rom(2231);
     when "100010111000" => data <= saw_rom(2232);
     when "100010111001" => data <= saw_rom(2233);
     when "100010111010" => data <= saw_rom(2234);
     when "100010111011" => data <= saw_rom(2235);
     when "100010111100" => data <= saw_rom(2236);
     when "100010111101" => data <= saw_rom(2237);
     when "100010111110" => data <= saw_rom(2238);
     when "100010111111" => data <= saw_rom(2239);
     when "100011000000" => data <= saw_rom(2240);
     when "100011000001" => data <= saw_rom(2241);
     when "100011000010" => data <= saw_rom(2242);
     when "100011000011" => data <= saw_rom(2243);
     when "100011000100" => data <= saw_rom(2244);
     when "100011000101" => data <= saw_rom(2245);
     when "100011000110" => data <= saw_rom(2246);
     when "100011000111" => data <= saw_rom(2247);
     when "100011001000" => data <= saw_rom(2248);
     when "100011001001" => data <= saw_rom(2249);
     when "100011001010" => data <= saw_rom(2250);
     when "100011001011" => data <= saw_rom(2251);
     when "100011001100" => data <= saw_rom(2252);
     when "100011001101" => data <= saw_rom(2253);
     when "100011001110" => data <= saw_rom(2254);
     when "100011001111" => data <= saw_rom(2255);
     when "100011010000" => data <= saw_rom(2256);
     when "100011010001" => data <= saw_rom(2257);
     when "100011010010" => data <= saw_rom(2258);
     when "100011010011" => data <= saw_rom(2259);
     when "100011010100" => data <= saw_rom(2260);
     when "100011010101" => data <= saw_rom(2261);
     when "100011010110" => data <= saw_rom(2262);
     when "100011010111" => data <= saw_rom(2263);
     when "100011011000" => data <= saw_rom(2264);
     when "100011011001" => data <= saw_rom(2265);
     when "100011011010" => data <= saw_rom(2266);
     when "100011011011" => data <= saw_rom(2267);
     when "100011011100" => data <= saw_rom(2268);
     when "100011011101" => data <= saw_rom(2269);
     when "100011011110" => data <= saw_rom(2270);
     when "100011011111" => data <= saw_rom(2271);
     when "100011100000" => data <= saw_rom(2272);
     when "100011100001" => data <= saw_rom(2273);
     when "100011100010" => data <= saw_rom(2274);
     when "100011100011" => data <= saw_rom(2275);
     when "100011100100" => data <= saw_rom(2276);
     when "100011100101" => data <= saw_rom(2277);
     when "100011100110" => data <= saw_rom(2278);
     when "100011100111" => data <= saw_rom(2279);
     when "100011101000" => data <= saw_rom(2280);
     when "100011101001" => data <= saw_rom(2281);
     when "100011101010" => data <= saw_rom(2282);
     when "100011101011" => data <= saw_rom(2283);
     when "100011101100" => data <= saw_rom(2284);
     when "100011101101" => data <= saw_rom(2285);
     when "100011101110" => data <= saw_rom(2286);
     when "100011101111" => data <= saw_rom(2287);
     when "100011110000" => data <= saw_rom(2288);
     when "100011110001" => data <= saw_rom(2289);
     when "100011110010" => data <= saw_rom(2290);
     when "100011110011" => data <= saw_rom(2291);
     when "100011110100" => data <= saw_rom(2292);
     when "100011110101" => data <= saw_rom(2293);
     when "100011110110" => data <= saw_rom(2294);
     when "100011110111" => data <= saw_rom(2295);
     when "100011111000" => data <= saw_rom(2296);
     when "100011111001" => data <= saw_rom(2297);
     when "100011111010" => data <= saw_rom(2298);
     when "100011111011" => data <= saw_rom(2299);
     when "100011111100" => data <= saw_rom(2300);
     when "100011111101" => data <= saw_rom(2301);
     when "100011111110" => data <= saw_rom(2302);
     when "100011111111" => data <= saw_rom(2303);
     when "100100000000" => data <= saw_rom(2304);
     when "100100000001" => data <= saw_rom(2305);
     when "100100000010" => data <= saw_rom(2306);
     when "100100000011" => data <= saw_rom(2307);
     when "100100000100" => data <= saw_rom(2308);
     when "100100000101" => data <= saw_rom(2309);
     when "100100000110" => data <= saw_rom(2310);
     when "100100000111" => data <= saw_rom(2311);
     when "100100001000" => data <= saw_rom(2312);
     when "100100001001" => data <= saw_rom(2313);
     when "100100001010" => data <= saw_rom(2314);
     when "100100001011" => data <= saw_rom(2315);
     when "100100001100" => data <= saw_rom(2316);
     when "100100001101" => data <= saw_rom(2317);
     when "100100001110" => data <= saw_rom(2318);
     when "100100001111" => data <= saw_rom(2319);
     when "100100010000" => data <= saw_rom(2320);
     when "100100010001" => data <= saw_rom(2321);
     when "100100010010" => data <= saw_rom(2322);
     when "100100010011" => data <= saw_rom(2323);
     when "100100010100" => data <= saw_rom(2324);
     when "100100010101" => data <= saw_rom(2325);
     when "100100010110" => data <= saw_rom(2326);
     when "100100010111" => data <= saw_rom(2327);
     when "100100011000" => data <= saw_rom(2328);
     when "100100011001" => data <= saw_rom(2329);
     when "100100011010" => data <= saw_rom(2330);
     when "100100011011" => data <= saw_rom(2331);
     when "100100011100" => data <= saw_rom(2332);
     when "100100011101" => data <= saw_rom(2333);
     when "100100011110" => data <= saw_rom(2334);
     when "100100011111" => data <= saw_rom(2335);
     when "100100100000" => data <= saw_rom(2336);
     when "100100100001" => data <= saw_rom(2337);
     when "100100100010" => data <= saw_rom(2338);
     when "100100100011" => data <= saw_rom(2339);
     when "100100100100" => data <= saw_rom(2340);
     when "100100100101" => data <= saw_rom(2341);
     when "100100100110" => data <= saw_rom(2342);
     when "100100100111" => data <= saw_rom(2343);
     when "100100101000" => data <= saw_rom(2344);
     when "100100101001" => data <= saw_rom(2345);
     when "100100101010" => data <= saw_rom(2346);
     when "100100101011" => data <= saw_rom(2347);
     when "100100101100" => data <= saw_rom(2348);
     when "100100101101" => data <= saw_rom(2349);
     when "100100101110" => data <= saw_rom(2350);
     when "100100101111" => data <= saw_rom(2351);
     when "100100110000" => data <= saw_rom(2352);
     when "100100110001" => data <= saw_rom(2353);
     when "100100110010" => data <= saw_rom(2354);
     when "100100110011" => data <= saw_rom(2355);
     when "100100110100" => data <= saw_rom(2356);
     when "100100110101" => data <= saw_rom(2357);
     when "100100110110" => data <= saw_rom(2358);
     when "100100110111" => data <= saw_rom(2359);
     when "100100111000" => data <= saw_rom(2360);
     when "100100111001" => data <= saw_rom(2361);
     when "100100111010" => data <= saw_rom(2362);
     when "100100111011" => data <= saw_rom(2363);
     when "100100111100" => data <= saw_rom(2364);
     when "100100111101" => data <= saw_rom(2365);
     when "100100111110" => data <= saw_rom(2366);
     when "100100111111" => data <= saw_rom(2367);
     when "100101000000" => data <= saw_rom(2368);
     when "100101000001" => data <= saw_rom(2369);
     when "100101000010" => data <= saw_rom(2370);
     when "100101000011" => data <= saw_rom(2371);
     when "100101000100" => data <= saw_rom(2372);
     when "100101000101" => data <= saw_rom(2373);
     when "100101000110" => data <= saw_rom(2374);
     when "100101000111" => data <= saw_rom(2375);
     when "100101001000" => data <= saw_rom(2376);
     when "100101001001" => data <= saw_rom(2377);
     when "100101001010" => data <= saw_rom(2378);
     when "100101001011" => data <= saw_rom(2379);
     when "100101001100" => data <= saw_rom(2380);
     when "100101001101" => data <= saw_rom(2381);
     when "100101001110" => data <= saw_rom(2382);
     when "100101001111" => data <= saw_rom(2383);
     when "100101010000" => data <= saw_rom(2384);
     when "100101010001" => data <= saw_rom(2385);
     when "100101010010" => data <= saw_rom(2386);
     when "100101010011" => data <= saw_rom(2387);
     when "100101010100" => data <= saw_rom(2388);
     when "100101010101" => data <= saw_rom(2389);
     when "100101010110" => data <= saw_rom(2390);
     when "100101010111" => data <= saw_rom(2391);
     when "100101011000" => data <= saw_rom(2392);
     when "100101011001" => data <= saw_rom(2393);
     when "100101011010" => data <= saw_rom(2394);
     when "100101011011" => data <= saw_rom(2395);
     when "100101011100" => data <= saw_rom(2396);
     when "100101011101" => data <= saw_rom(2397);
     when "100101011110" => data <= saw_rom(2398);
     when "100101011111" => data <= saw_rom(2399);
     when "100101100000" => data <= saw_rom(2400);
     when "100101100001" => data <= saw_rom(2401);
     when "100101100010" => data <= saw_rom(2402);
     when "100101100011" => data <= saw_rom(2403);
     when "100101100100" => data <= saw_rom(2404);
     when "100101100101" => data <= saw_rom(2405);
     when "100101100110" => data <= saw_rom(2406);
     when "100101100111" => data <= saw_rom(2407);
     when "100101101000" => data <= saw_rom(2408);
     when "100101101001" => data <= saw_rom(2409);
     when "100101101010" => data <= saw_rom(2410);
     when "100101101011" => data <= saw_rom(2411);
     when "100101101100" => data <= saw_rom(2412);
     when "100101101101" => data <= saw_rom(2413);
     when "100101101110" => data <= saw_rom(2414);
     when "100101101111" => data <= saw_rom(2415);
     when "100101110000" => data <= saw_rom(2416);
     when "100101110001" => data <= saw_rom(2417);
     when "100101110010" => data <= saw_rom(2418);
     when "100101110011" => data <= saw_rom(2419);
     when "100101110100" => data <= saw_rom(2420);
     when "100101110101" => data <= saw_rom(2421);
     when "100101110110" => data <= saw_rom(2422);
     when "100101110111" => data <= saw_rom(2423);
     when "100101111000" => data <= saw_rom(2424);
     when "100101111001" => data <= saw_rom(2425);
     when "100101111010" => data <= saw_rom(2426);
     when "100101111011" => data <= saw_rom(2427);
     when "100101111100" => data <= saw_rom(2428);
     when "100101111101" => data <= saw_rom(2429);
     when "100101111110" => data <= saw_rom(2430);
     when "100101111111" => data <= saw_rom(2431);
     when "100110000000" => data <= saw_rom(2432);
     when "100110000001" => data <= saw_rom(2433);
     when "100110000010" => data <= saw_rom(2434);
     when "100110000011" => data <= saw_rom(2435);
     when "100110000100" => data <= saw_rom(2436);
     when "100110000101" => data <= saw_rom(2437);
     when "100110000110" => data <= saw_rom(2438);
     when "100110000111" => data <= saw_rom(2439);
     when "100110001000" => data <= saw_rom(2440);
     when "100110001001" => data <= saw_rom(2441);
     when "100110001010" => data <= saw_rom(2442);
     when "100110001011" => data <= saw_rom(2443);
     when "100110001100" => data <= saw_rom(2444);
     when "100110001101" => data <= saw_rom(2445);
     when "100110001110" => data <= saw_rom(2446);
     when "100110001111" => data <= saw_rom(2447);
     when "100110010000" => data <= saw_rom(2448);
     when "100110010001" => data <= saw_rom(2449);
     when "100110010010" => data <= saw_rom(2450);
     when "100110010011" => data <= saw_rom(2451);
     when "100110010100" => data <= saw_rom(2452);
     when "100110010101" => data <= saw_rom(2453);
     when "100110010110" => data <= saw_rom(2454);
     when "100110010111" => data <= saw_rom(2455);
     when "100110011000" => data <= saw_rom(2456);
     when "100110011001" => data <= saw_rom(2457);
     when "100110011010" => data <= saw_rom(2458);
     when "100110011011" => data <= saw_rom(2459);
     when "100110011100" => data <= saw_rom(2460);
     when "100110011101" => data <= saw_rom(2461);
     when "100110011110" => data <= saw_rom(2462);
     when "100110011111" => data <= saw_rom(2463);
     when "100110100000" => data <= saw_rom(2464);
     when "100110100001" => data <= saw_rom(2465);
     when "100110100010" => data <= saw_rom(2466);
     when "100110100011" => data <= saw_rom(2467);
     when "100110100100" => data <= saw_rom(2468);
     when "100110100101" => data <= saw_rom(2469);
     when "100110100110" => data <= saw_rom(2470);
     when "100110100111" => data <= saw_rom(2471);
     when "100110101000" => data <= saw_rom(2472);
     when "100110101001" => data <= saw_rom(2473);
     when "100110101010" => data <= saw_rom(2474);
     when "100110101011" => data <= saw_rom(2475);
     when "100110101100" => data <= saw_rom(2476);
     when "100110101101" => data <= saw_rom(2477);
     when "100110101110" => data <= saw_rom(2478);
     when "100110101111" => data <= saw_rom(2479);
     when "100110110000" => data <= saw_rom(2480);
     when "100110110001" => data <= saw_rom(2481);
     when "100110110010" => data <= saw_rom(2482);
     when "100110110011" => data <= saw_rom(2483);
     when "100110110100" => data <= saw_rom(2484);
     when "100110110101" => data <= saw_rom(2485);
     when "100110110110" => data <= saw_rom(2486);
     when "100110110111" => data <= saw_rom(2487);
     when "100110111000" => data <= saw_rom(2488);
     when "100110111001" => data <= saw_rom(2489);
     when "100110111010" => data <= saw_rom(2490);
     when "100110111011" => data <= saw_rom(2491);
     when "100110111100" => data <= saw_rom(2492);
     when "100110111101" => data <= saw_rom(2493);
     when "100110111110" => data <= saw_rom(2494);
     when "100110111111" => data <= saw_rom(2495);
     when "100111000000" => data <= saw_rom(2496);
     when "100111000001" => data <= saw_rom(2497);
     when "100111000010" => data <= saw_rom(2498);
     when "100111000011" => data <= saw_rom(2499);
     when "100111000100" => data <= saw_rom(2500);
     when "100111000101" => data <= saw_rom(2501);
     when "100111000110" => data <= saw_rom(2502);
     when "100111000111" => data <= saw_rom(2503);
     when "100111001000" => data <= saw_rom(2504);
     when "100111001001" => data <= saw_rom(2505);
     when "100111001010" => data <= saw_rom(2506);
     when "100111001011" => data <= saw_rom(2507);
     when "100111001100" => data <= saw_rom(2508);
     when "100111001101" => data <= saw_rom(2509);
     when "100111001110" => data <= saw_rom(2510);
     when "100111001111" => data <= saw_rom(2511);
     when "100111010000" => data <= saw_rom(2512);
     when "100111010001" => data <= saw_rom(2513);
     when "100111010010" => data <= saw_rom(2514);
     when "100111010011" => data <= saw_rom(2515);
     when "100111010100" => data <= saw_rom(2516);
     when "100111010101" => data <= saw_rom(2517);
     when "100111010110" => data <= saw_rom(2518);
     when "100111010111" => data <= saw_rom(2519);
     when "100111011000" => data <= saw_rom(2520);
     when "100111011001" => data <= saw_rom(2521);
     when "100111011010" => data <= saw_rom(2522);
     when "100111011011" => data <= saw_rom(2523);
     when "100111011100" => data <= saw_rom(2524);
     when "100111011101" => data <= saw_rom(2525);
     when "100111011110" => data <= saw_rom(2526);
     when "100111011111" => data <= saw_rom(2527);
     when "100111100000" => data <= saw_rom(2528);
     when "100111100001" => data <= saw_rom(2529);
     when "100111100010" => data <= saw_rom(2530);
     when "100111100011" => data <= saw_rom(2531);
     when "100111100100" => data <= saw_rom(2532);
     when "100111100101" => data <= saw_rom(2533);
     when "100111100110" => data <= saw_rom(2534);
     when "100111100111" => data <= saw_rom(2535);
     when "100111101000" => data <= saw_rom(2536);
     when "100111101001" => data <= saw_rom(2537);
     when "100111101010" => data <= saw_rom(2538);
     when "100111101011" => data <= saw_rom(2539);
     when "100111101100" => data <= saw_rom(2540);
     when "100111101101" => data <= saw_rom(2541);
     when "100111101110" => data <= saw_rom(2542);
     when "100111101111" => data <= saw_rom(2543);
     when "100111110000" => data <= saw_rom(2544);
     when "100111110001" => data <= saw_rom(2545);
     when "100111110010" => data <= saw_rom(2546);
     when "100111110011" => data <= saw_rom(2547);
     when "100111110100" => data <= saw_rom(2548);
     when "100111110101" => data <= saw_rom(2549);
     when "100111110110" => data <= saw_rom(2550);
     when "100111110111" => data <= saw_rom(2551);
     when "100111111000" => data <= saw_rom(2552);
     when "100111111001" => data <= saw_rom(2553);
     when "100111111010" => data <= saw_rom(2554);
     when "100111111011" => data <= saw_rom(2555);
     when "100111111100" => data <= saw_rom(2556);
     when "100111111101" => data <= saw_rom(2557);
     when "100111111110" => data <= saw_rom(2558);
     when "100111111111" => data <= saw_rom(2559);
     when "101000000000" => data <= saw_rom(2560);
     when "101000000001" => data <= saw_rom(2561);
     when "101000000010" => data <= saw_rom(2562);
     when "101000000011" => data <= saw_rom(2563);
     when "101000000100" => data <= saw_rom(2564);
     when "101000000101" => data <= saw_rom(2565);
     when "101000000110" => data <= saw_rom(2566);
     when "101000000111" => data <= saw_rom(2567);
     when "101000001000" => data <= saw_rom(2568);
     when "101000001001" => data <= saw_rom(2569);
     when "101000001010" => data <= saw_rom(2570);
     when "101000001011" => data <= saw_rom(2571);
     when "101000001100" => data <= saw_rom(2572);
     when "101000001101" => data <= saw_rom(2573);
     when "101000001110" => data <= saw_rom(2574);
     when "101000001111" => data <= saw_rom(2575);
     when "101000010000" => data <= saw_rom(2576);
     when "101000010001" => data <= saw_rom(2577);
     when "101000010010" => data <= saw_rom(2578);
     when "101000010011" => data <= saw_rom(2579);
     when "101000010100" => data <= saw_rom(2580);
     when "101000010101" => data <= saw_rom(2581);
     when "101000010110" => data <= saw_rom(2582);
     when "101000010111" => data <= saw_rom(2583);
     when "101000011000" => data <= saw_rom(2584);
     when "101000011001" => data <= saw_rom(2585);
     when "101000011010" => data <= saw_rom(2586);
     when "101000011011" => data <= saw_rom(2587);
     when "101000011100" => data <= saw_rom(2588);
     when "101000011101" => data <= saw_rom(2589);
     when "101000011110" => data <= saw_rom(2590);
     when "101000011111" => data <= saw_rom(2591);
     when "101000100000" => data <= saw_rom(2592);
     when "101000100001" => data <= saw_rom(2593);
     when "101000100010" => data <= saw_rom(2594);
     when "101000100011" => data <= saw_rom(2595);
     when "101000100100" => data <= saw_rom(2596);
     when "101000100101" => data <= saw_rom(2597);
     when "101000100110" => data <= saw_rom(2598);
     when "101000100111" => data <= saw_rom(2599);
     when "101000101000" => data <= saw_rom(2600);
     when "101000101001" => data <= saw_rom(2601);
     when "101000101010" => data <= saw_rom(2602);
     when "101000101011" => data <= saw_rom(2603);
     when "101000101100" => data <= saw_rom(2604);
     when "101000101101" => data <= saw_rom(2605);
     when "101000101110" => data <= saw_rom(2606);
     when "101000101111" => data <= saw_rom(2607);
     when "101000110000" => data <= saw_rom(2608);
     when "101000110001" => data <= saw_rom(2609);
     when "101000110010" => data <= saw_rom(2610);
     when "101000110011" => data <= saw_rom(2611);
     when "101000110100" => data <= saw_rom(2612);
     when "101000110101" => data <= saw_rom(2613);
     when "101000110110" => data <= saw_rom(2614);
     when "101000110111" => data <= saw_rom(2615);
     when "101000111000" => data <= saw_rom(2616);
     when "101000111001" => data <= saw_rom(2617);
     when "101000111010" => data <= saw_rom(2618);
     when "101000111011" => data <= saw_rom(2619);
     when "101000111100" => data <= saw_rom(2620);
     when "101000111101" => data <= saw_rom(2621);
     when "101000111110" => data <= saw_rom(2622);
     when "101000111111" => data <= saw_rom(2623);
     when "101001000000" => data <= saw_rom(2624);
     when "101001000001" => data <= saw_rom(2625);
     when "101001000010" => data <= saw_rom(2626);
     when "101001000011" => data <= saw_rom(2627);
     when "101001000100" => data <= saw_rom(2628);
     when "101001000101" => data <= saw_rom(2629);
     when "101001000110" => data <= saw_rom(2630);
     when "101001000111" => data <= saw_rom(2631);
     when "101001001000" => data <= saw_rom(2632);
     when "101001001001" => data <= saw_rom(2633);
     when "101001001010" => data <= saw_rom(2634);
     when "101001001011" => data <= saw_rom(2635);
     when "101001001100" => data <= saw_rom(2636);
     when "101001001101" => data <= saw_rom(2637);
     when "101001001110" => data <= saw_rom(2638);
     when "101001001111" => data <= saw_rom(2639);
     when "101001010000" => data <= saw_rom(2640);
     when "101001010001" => data <= saw_rom(2641);
     when "101001010010" => data <= saw_rom(2642);
     when "101001010011" => data <= saw_rom(2643);
     when "101001010100" => data <= saw_rom(2644);
     when "101001010101" => data <= saw_rom(2645);
     when "101001010110" => data <= saw_rom(2646);
     when "101001010111" => data <= saw_rom(2647);
     when "101001011000" => data <= saw_rom(2648);
     when "101001011001" => data <= saw_rom(2649);
     when "101001011010" => data <= saw_rom(2650);
     when "101001011011" => data <= saw_rom(2651);
     when "101001011100" => data <= saw_rom(2652);
     when "101001011101" => data <= saw_rom(2653);
     when "101001011110" => data <= saw_rom(2654);
     when "101001011111" => data <= saw_rom(2655);
     when "101001100000" => data <= saw_rom(2656);
     when "101001100001" => data <= saw_rom(2657);
     when "101001100010" => data <= saw_rom(2658);
     when "101001100011" => data <= saw_rom(2659);
     when "101001100100" => data <= saw_rom(2660);
     when "101001100101" => data <= saw_rom(2661);
     when "101001100110" => data <= saw_rom(2662);
     when "101001100111" => data <= saw_rom(2663);
     when "101001101000" => data <= saw_rom(2664);
     when "101001101001" => data <= saw_rom(2665);
     when "101001101010" => data <= saw_rom(2666);
     when "101001101011" => data <= saw_rom(2667);
     when "101001101100" => data <= saw_rom(2668);
     when "101001101101" => data <= saw_rom(2669);
     when "101001101110" => data <= saw_rom(2670);
     when "101001101111" => data <= saw_rom(2671);
     when "101001110000" => data <= saw_rom(2672);
     when "101001110001" => data <= saw_rom(2673);
     when "101001110010" => data <= saw_rom(2674);
     when "101001110011" => data <= saw_rom(2675);
     when "101001110100" => data <= saw_rom(2676);
     when "101001110101" => data <= saw_rom(2677);
     when "101001110110" => data <= saw_rom(2678);
     when "101001110111" => data <= saw_rom(2679);
     when "101001111000" => data <= saw_rom(2680);
     when "101001111001" => data <= saw_rom(2681);
     when "101001111010" => data <= saw_rom(2682);
     when "101001111011" => data <= saw_rom(2683);
     when "101001111100" => data <= saw_rom(2684);
     when "101001111101" => data <= saw_rom(2685);
     when "101001111110" => data <= saw_rom(2686);
     when "101001111111" => data <= saw_rom(2687);
     when "101010000000" => data <= saw_rom(2688);
     when "101010000001" => data <= saw_rom(2689);
     when "101010000010" => data <= saw_rom(2690);
     when "101010000011" => data <= saw_rom(2691);
     when "101010000100" => data <= saw_rom(2692);
     when "101010000101" => data <= saw_rom(2693);
     when "101010000110" => data <= saw_rom(2694);
     when "101010000111" => data <= saw_rom(2695);
     when "101010001000" => data <= saw_rom(2696);
     when "101010001001" => data <= saw_rom(2697);
     when "101010001010" => data <= saw_rom(2698);
     when "101010001011" => data <= saw_rom(2699);
     when "101010001100" => data <= saw_rom(2700);
     when "101010001101" => data <= saw_rom(2701);
     when "101010001110" => data <= saw_rom(2702);
     when "101010001111" => data <= saw_rom(2703);
     when "101010010000" => data <= saw_rom(2704);
     when "101010010001" => data <= saw_rom(2705);
     when "101010010010" => data <= saw_rom(2706);
     when "101010010011" => data <= saw_rom(2707);
     when "101010010100" => data <= saw_rom(2708);
     when "101010010101" => data <= saw_rom(2709);
     when "101010010110" => data <= saw_rom(2710);
     when "101010010111" => data <= saw_rom(2711);
     when "101010011000" => data <= saw_rom(2712);
     when "101010011001" => data <= saw_rom(2713);
     when "101010011010" => data <= saw_rom(2714);
     when "101010011011" => data <= saw_rom(2715);
     when "101010011100" => data <= saw_rom(2716);
     when "101010011101" => data <= saw_rom(2717);
     when "101010011110" => data <= saw_rom(2718);
     when "101010011111" => data <= saw_rom(2719);
     when "101010100000" => data <= saw_rom(2720);
     when "101010100001" => data <= saw_rom(2721);
     when "101010100010" => data <= saw_rom(2722);
     when "101010100011" => data <= saw_rom(2723);
     when "101010100100" => data <= saw_rom(2724);
     when "101010100101" => data <= saw_rom(2725);
     when "101010100110" => data <= saw_rom(2726);
     when "101010100111" => data <= saw_rom(2727);
     when "101010101000" => data <= saw_rom(2728);
     when "101010101001" => data <= saw_rom(2729);
     when "101010101010" => data <= saw_rom(2730);
     when "101010101011" => data <= saw_rom(2731);
     when "101010101100" => data <= saw_rom(2732);
     when "101010101101" => data <= saw_rom(2733);
     when "101010101110" => data <= saw_rom(2734);
     when "101010101111" => data <= saw_rom(2735);
     when "101010110000" => data <= saw_rom(2736);
     when "101010110001" => data <= saw_rom(2737);
     when "101010110010" => data <= saw_rom(2738);
     when "101010110011" => data <= saw_rom(2739);
     when "101010110100" => data <= saw_rom(2740);
     when "101010110101" => data <= saw_rom(2741);
     when "101010110110" => data <= saw_rom(2742);
     when "101010110111" => data <= saw_rom(2743);
     when "101010111000" => data <= saw_rom(2744);
     when "101010111001" => data <= saw_rom(2745);
     when "101010111010" => data <= saw_rom(2746);
     when "101010111011" => data <= saw_rom(2747);
     when "101010111100" => data <= saw_rom(2748);
     when "101010111101" => data <= saw_rom(2749);
     when "101010111110" => data <= saw_rom(2750);
     when "101010111111" => data <= saw_rom(2751);
     when "101011000000" => data <= saw_rom(2752);
     when "101011000001" => data <= saw_rom(2753);
     when "101011000010" => data <= saw_rom(2754);
     when "101011000011" => data <= saw_rom(2755);
     when "101011000100" => data <= saw_rom(2756);
     when "101011000101" => data <= saw_rom(2757);
     when "101011000110" => data <= saw_rom(2758);
     when "101011000111" => data <= saw_rom(2759);
     when "101011001000" => data <= saw_rom(2760);
     when "101011001001" => data <= saw_rom(2761);
     when "101011001010" => data <= saw_rom(2762);
     when "101011001011" => data <= saw_rom(2763);
     when "101011001100" => data <= saw_rom(2764);
     when "101011001101" => data <= saw_rom(2765);
     when "101011001110" => data <= saw_rom(2766);
     when "101011001111" => data <= saw_rom(2767);
     when "101011010000" => data <= saw_rom(2768);
     when "101011010001" => data <= saw_rom(2769);
     when "101011010010" => data <= saw_rom(2770);
     when "101011010011" => data <= saw_rom(2771);
     when "101011010100" => data <= saw_rom(2772);
     when "101011010101" => data <= saw_rom(2773);
     when "101011010110" => data <= saw_rom(2774);
     when "101011010111" => data <= saw_rom(2775);
     when "101011011000" => data <= saw_rom(2776);
     when "101011011001" => data <= saw_rom(2777);
     when "101011011010" => data <= saw_rom(2778);
     when "101011011011" => data <= saw_rom(2779);
     when "101011011100" => data <= saw_rom(2780);
     when "101011011101" => data <= saw_rom(2781);
     when "101011011110" => data <= saw_rom(2782);
     when "101011011111" => data <= saw_rom(2783);
     when "101011100000" => data <= saw_rom(2784);
     when "101011100001" => data <= saw_rom(2785);
     when "101011100010" => data <= saw_rom(2786);
     when "101011100011" => data <= saw_rom(2787);
     when "101011100100" => data <= saw_rom(2788);
     when "101011100101" => data <= saw_rom(2789);
     when "101011100110" => data <= saw_rom(2790);
     when "101011100111" => data <= saw_rom(2791);
     when "101011101000" => data <= saw_rom(2792);
     when "101011101001" => data <= saw_rom(2793);
     when "101011101010" => data <= saw_rom(2794);
     when "101011101011" => data <= saw_rom(2795);
     when "101011101100" => data <= saw_rom(2796);
     when "101011101101" => data <= saw_rom(2797);
     when "101011101110" => data <= saw_rom(2798);
     when "101011101111" => data <= saw_rom(2799);
     when "101011110000" => data <= saw_rom(2800);
     when "101011110001" => data <= saw_rom(2801);
     when "101011110010" => data <= saw_rom(2802);
     when "101011110011" => data <= saw_rom(2803);
     when "101011110100" => data <= saw_rom(2804);
     when "101011110101" => data <= saw_rom(2805);
     when "101011110110" => data <= saw_rom(2806);
     when "101011110111" => data <= saw_rom(2807);
     when "101011111000" => data <= saw_rom(2808);
     when "101011111001" => data <= saw_rom(2809);
     when "101011111010" => data <= saw_rom(2810);
     when "101011111011" => data <= saw_rom(2811);
     when "101011111100" => data <= saw_rom(2812);
     when "101011111101" => data <= saw_rom(2813);
     when "101011111110" => data <= saw_rom(2814);
     when "101011111111" => data <= saw_rom(2815);
     when "101100000000" => data <= saw_rom(2816);
     when "101100000001" => data <= saw_rom(2817);
     when "101100000010" => data <= saw_rom(2818);
     when "101100000011" => data <= saw_rom(2819);
     when "101100000100" => data <= saw_rom(2820);
     when "101100000101" => data <= saw_rom(2821);
     when "101100000110" => data <= saw_rom(2822);
     when "101100000111" => data <= saw_rom(2823);
     when "101100001000" => data <= saw_rom(2824);
     when "101100001001" => data <= saw_rom(2825);
     when "101100001010" => data <= saw_rom(2826);
     when "101100001011" => data <= saw_rom(2827);
     when "101100001100" => data <= saw_rom(2828);
     when "101100001101" => data <= saw_rom(2829);
     when "101100001110" => data <= saw_rom(2830);
     when "101100001111" => data <= saw_rom(2831);
     when "101100010000" => data <= saw_rom(2832);
     when "101100010001" => data <= saw_rom(2833);
     when "101100010010" => data <= saw_rom(2834);
     when "101100010011" => data <= saw_rom(2835);
     when "101100010100" => data <= saw_rom(2836);
     when "101100010101" => data <= saw_rom(2837);
     when "101100010110" => data <= saw_rom(2838);
     when "101100010111" => data <= saw_rom(2839);
     when "101100011000" => data <= saw_rom(2840);
     when "101100011001" => data <= saw_rom(2841);
     when "101100011010" => data <= saw_rom(2842);
     when "101100011011" => data <= saw_rom(2843);
     when "101100011100" => data <= saw_rom(2844);
     when "101100011101" => data <= saw_rom(2845);
     when "101100011110" => data <= saw_rom(2846);
     when "101100011111" => data <= saw_rom(2847);
     when "101100100000" => data <= saw_rom(2848);
     when "101100100001" => data <= saw_rom(2849);
     when "101100100010" => data <= saw_rom(2850);
     when "101100100011" => data <= saw_rom(2851);
     when "101100100100" => data <= saw_rom(2852);
     when "101100100101" => data <= saw_rom(2853);
     when "101100100110" => data <= saw_rom(2854);
     when "101100100111" => data <= saw_rom(2855);
     when "101100101000" => data <= saw_rom(2856);
     when "101100101001" => data <= saw_rom(2857);
     when "101100101010" => data <= saw_rom(2858);
     when "101100101011" => data <= saw_rom(2859);
     when "101100101100" => data <= saw_rom(2860);
     when "101100101101" => data <= saw_rom(2861);
     when "101100101110" => data <= saw_rom(2862);
     when "101100101111" => data <= saw_rom(2863);
     when "101100110000" => data <= saw_rom(2864);
     when "101100110001" => data <= saw_rom(2865);
     when "101100110010" => data <= saw_rom(2866);
     when "101100110011" => data <= saw_rom(2867);
     when "101100110100" => data <= saw_rom(2868);
     when "101100110101" => data <= saw_rom(2869);
     when "101100110110" => data <= saw_rom(2870);
     when "101100110111" => data <= saw_rom(2871);
     when "101100111000" => data <= saw_rom(2872);
     when "101100111001" => data <= saw_rom(2873);
     when "101100111010" => data <= saw_rom(2874);
     when "101100111011" => data <= saw_rom(2875);
     when "101100111100" => data <= saw_rom(2876);
     when "101100111101" => data <= saw_rom(2877);
     when "101100111110" => data <= saw_rom(2878);
     when "101100111111" => data <= saw_rom(2879);
     when "101101000000" => data <= saw_rom(2880);
     when "101101000001" => data <= saw_rom(2881);
     when "101101000010" => data <= saw_rom(2882);
     when "101101000011" => data <= saw_rom(2883);
     when "101101000100" => data <= saw_rom(2884);
     when "101101000101" => data <= saw_rom(2885);
     when "101101000110" => data <= saw_rom(2886);
     when "101101000111" => data <= saw_rom(2887);
     when "101101001000" => data <= saw_rom(2888);
     when "101101001001" => data <= saw_rom(2889);
     when "101101001010" => data <= saw_rom(2890);
     when "101101001011" => data <= saw_rom(2891);
     when "101101001100" => data <= saw_rom(2892);
     when "101101001101" => data <= saw_rom(2893);
     when "101101001110" => data <= saw_rom(2894);
     when "101101001111" => data <= saw_rom(2895);
     when "101101010000" => data <= saw_rom(2896);
     when "101101010001" => data <= saw_rom(2897);
     when "101101010010" => data <= saw_rom(2898);
     when "101101010011" => data <= saw_rom(2899);
     when "101101010100" => data <= saw_rom(2900);
     when "101101010101" => data <= saw_rom(2901);
     when "101101010110" => data <= saw_rom(2902);
     when "101101010111" => data <= saw_rom(2903);
     when "101101011000" => data <= saw_rom(2904);
     when "101101011001" => data <= saw_rom(2905);
     when "101101011010" => data <= saw_rom(2906);
     when "101101011011" => data <= saw_rom(2907);
     when "101101011100" => data <= saw_rom(2908);
     when "101101011101" => data <= saw_rom(2909);
     when "101101011110" => data <= saw_rom(2910);
     when "101101011111" => data <= saw_rom(2911);
     when "101101100000" => data <= saw_rom(2912);
     when "101101100001" => data <= saw_rom(2913);
     when "101101100010" => data <= saw_rom(2914);
     when "101101100011" => data <= saw_rom(2915);
     when "101101100100" => data <= saw_rom(2916);
     when "101101100101" => data <= saw_rom(2917);
     when "101101100110" => data <= saw_rom(2918);
     when "101101100111" => data <= saw_rom(2919);
     when "101101101000" => data <= saw_rom(2920);
     when "101101101001" => data <= saw_rom(2921);
     when "101101101010" => data <= saw_rom(2922);
     when "101101101011" => data <= saw_rom(2923);
     when "101101101100" => data <= saw_rom(2924);
     when "101101101101" => data <= saw_rom(2925);
     when "101101101110" => data <= saw_rom(2926);
     when "101101101111" => data <= saw_rom(2927);
     when "101101110000" => data <= saw_rom(2928);
     when "101101110001" => data <= saw_rom(2929);
     when "101101110010" => data <= saw_rom(2930);
     when "101101110011" => data <= saw_rom(2931);
     when "101101110100" => data <= saw_rom(2932);
     when "101101110101" => data <= saw_rom(2933);
     when "101101110110" => data <= saw_rom(2934);
     when "101101110111" => data <= saw_rom(2935);
     when "101101111000" => data <= saw_rom(2936);
     when "101101111001" => data <= saw_rom(2937);
     when "101101111010" => data <= saw_rom(2938);
     when "101101111011" => data <= saw_rom(2939);
     when "101101111100" => data <= saw_rom(2940);
     when "101101111101" => data <= saw_rom(2941);
     when "101101111110" => data <= saw_rom(2942);
     when "101101111111" => data <= saw_rom(2943);
     when "101110000000" => data <= saw_rom(2944);
     when "101110000001" => data <= saw_rom(2945);
     when "101110000010" => data <= saw_rom(2946);
     when "101110000011" => data <= saw_rom(2947);
     when "101110000100" => data <= saw_rom(2948);
     when "101110000101" => data <= saw_rom(2949);
     when "101110000110" => data <= saw_rom(2950);
     when "101110000111" => data <= saw_rom(2951);
     when "101110001000" => data <= saw_rom(2952);
     when "101110001001" => data <= saw_rom(2953);
     when "101110001010" => data <= saw_rom(2954);
     when "101110001011" => data <= saw_rom(2955);
     when "101110001100" => data <= saw_rom(2956);
     when "101110001101" => data <= saw_rom(2957);
     when "101110001110" => data <= saw_rom(2958);
     when "101110001111" => data <= saw_rom(2959);
     when "101110010000" => data <= saw_rom(2960);
     when "101110010001" => data <= saw_rom(2961);
     when "101110010010" => data <= saw_rom(2962);
     when "101110010011" => data <= saw_rom(2963);
     when "101110010100" => data <= saw_rom(2964);
     when "101110010101" => data <= saw_rom(2965);
     when "101110010110" => data <= saw_rom(2966);
     when "101110010111" => data <= saw_rom(2967);
     when "101110011000" => data <= saw_rom(2968);
     when "101110011001" => data <= saw_rom(2969);
     when "101110011010" => data <= saw_rom(2970);
     when "101110011011" => data <= saw_rom(2971);
     when "101110011100" => data <= saw_rom(2972);
     when "101110011101" => data <= saw_rom(2973);
     when "101110011110" => data <= saw_rom(2974);
     when "101110011111" => data <= saw_rom(2975);
     when "101110100000" => data <= saw_rom(2976);
     when "101110100001" => data <= saw_rom(2977);
     when "101110100010" => data <= saw_rom(2978);
     when "101110100011" => data <= saw_rom(2979);
     when "101110100100" => data <= saw_rom(2980);
     when "101110100101" => data <= saw_rom(2981);
     when "101110100110" => data <= saw_rom(2982);
     when "101110100111" => data <= saw_rom(2983);
     when "101110101000" => data <= saw_rom(2984);
     when "101110101001" => data <= saw_rom(2985);
     when "101110101010" => data <= saw_rom(2986);
     when "101110101011" => data <= saw_rom(2987);
     when "101110101100" => data <= saw_rom(2988);
     when "101110101101" => data <= saw_rom(2989);
     when "101110101110" => data <= saw_rom(2990);
     when "101110101111" => data <= saw_rom(2991);
     when "101110110000" => data <= saw_rom(2992);
     when "101110110001" => data <= saw_rom(2993);
     when "101110110010" => data <= saw_rom(2994);
     when "101110110011" => data <= saw_rom(2995);
     when "101110110100" => data <= saw_rom(2996);
     when "101110110101" => data <= saw_rom(2997);
     when "101110110110" => data <= saw_rom(2998);
     when "101110110111" => data <= saw_rom(2999);
     when "101110111000" => data <= saw_rom(3000);
     when "101110111001" => data <= saw_rom(3001);
     when "101110111010" => data <= saw_rom(3002);
     when "101110111011" => data <= saw_rom(3003);
     when "101110111100" => data <= saw_rom(3004);
     when "101110111101" => data <= saw_rom(3005);
     when "101110111110" => data <= saw_rom(3006);
     when "101110111111" => data <= saw_rom(3007);
     when "101111000000" => data <= saw_rom(3008);
     when "101111000001" => data <= saw_rom(3009);
     when "101111000010" => data <= saw_rom(3010);
     when "101111000011" => data <= saw_rom(3011);
     when "101111000100" => data <= saw_rom(3012);
     when "101111000101" => data <= saw_rom(3013);
     when "101111000110" => data <= saw_rom(3014);
     when "101111000111" => data <= saw_rom(3015);
     when "101111001000" => data <= saw_rom(3016);
     when "101111001001" => data <= saw_rom(3017);
     when "101111001010" => data <= saw_rom(3018);
     when "101111001011" => data <= saw_rom(3019);
     when "101111001100" => data <= saw_rom(3020);
     when "101111001101" => data <= saw_rom(3021);
     when "101111001110" => data <= saw_rom(3022);
     when "101111001111" => data <= saw_rom(3023);
     when "101111010000" => data <= saw_rom(3024);
     when "101111010001" => data <= saw_rom(3025);
     when "101111010010" => data <= saw_rom(3026);
     when "101111010011" => data <= saw_rom(3027);
     when "101111010100" => data <= saw_rom(3028);
     when "101111010101" => data <= saw_rom(3029);
     when "101111010110" => data <= saw_rom(3030);
     when "101111010111" => data <= saw_rom(3031);
     when "101111011000" => data <= saw_rom(3032);
     when "101111011001" => data <= saw_rom(3033);
     when "101111011010" => data <= saw_rom(3034);
     when "101111011011" => data <= saw_rom(3035);
     when "101111011100" => data <= saw_rom(3036);
     when "101111011101" => data <= saw_rom(3037);
     when "101111011110" => data <= saw_rom(3038);
     when "101111011111" => data <= saw_rom(3039);
     when "101111100000" => data <= saw_rom(3040);
     when "101111100001" => data <= saw_rom(3041);
     when "101111100010" => data <= saw_rom(3042);
     when "101111100011" => data <= saw_rom(3043);
     when "101111100100" => data <= saw_rom(3044);
     when "101111100101" => data <= saw_rom(3045);
     when "101111100110" => data <= saw_rom(3046);
     when "101111100111" => data <= saw_rom(3047);
     when "101111101000" => data <= saw_rom(3048);
     when "101111101001" => data <= saw_rom(3049);
     when "101111101010" => data <= saw_rom(3050);
     when "101111101011" => data <= saw_rom(3051);
     when "101111101100" => data <= saw_rom(3052);
     when "101111101101" => data <= saw_rom(3053);
     when "101111101110" => data <= saw_rom(3054);
     when "101111101111" => data <= saw_rom(3055);
     when "101111110000" => data <= saw_rom(3056);
     when "101111110001" => data <= saw_rom(3057);
     when "101111110010" => data <= saw_rom(3058);
     when "101111110011" => data <= saw_rom(3059);
     when "101111110100" => data <= saw_rom(3060);
     when "101111110101" => data <= saw_rom(3061);
     when "101111110110" => data <= saw_rom(3062);
     when "101111110111" => data <= saw_rom(3063);
     when "101111111000" => data <= saw_rom(3064);
     when "101111111001" => data <= saw_rom(3065);
     when "101111111010" => data <= saw_rom(3066);
     when "101111111011" => data <= saw_rom(3067);
     when "101111111100" => data <= saw_rom(3068);
     when "101111111101" => data <= saw_rom(3069);
     when "101111111110" => data <= saw_rom(3070);
     when "101111111111" => data <= saw_rom(3071);
     when "110000000000" => data <= saw_rom(3072);
     when "110000000001" => data <= saw_rom(3073);
     when "110000000010" => data <= saw_rom(3074);
     when "110000000011" => data <= saw_rom(3075);
     when "110000000100" => data <= saw_rom(3076);
     when "110000000101" => data <= saw_rom(3077);
     when "110000000110" => data <= saw_rom(3078);
     when "110000000111" => data <= saw_rom(3079);
     when "110000001000" => data <= saw_rom(3080);
     when "110000001001" => data <= saw_rom(3081);
     when "110000001010" => data <= saw_rom(3082);
     when "110000001011" => data <= saw_rom(3083);
     when "110000001100" => data <= saw_rom(3084);
     when "110000001101" => data <= saw_rom(3085);
     when "110000001110" => data <= saw_rom(3086);
     when "110000001111" => data <= saw_rom(3087);
     when "110000010000" => data <= saw_rom(3088);
     when "110000010001" => data <= saw_rom(3089);
     when "110000010010" => data <= saw_rom(3090);
     when "110000010011" => data <= saw_rom(3091);
     when "110000010100" => data <= saw_rom(3092);
     when "110000010101" => data <= saw_rom(3093);
     when "110000010110" => data <= saw_rom(3094);
     when "110000010111" => data <= saw_rom(3095);
     when "110000011000" => data <= saw_rom(3096);
     when "110000011001" => data <= saw_rom(3097);
     when "110000011010" => data <= saw_rom(3098);
     when "110000011011" => data <= saw_rom(3099);
     when "110000011100" => data <= saw_rom(3100);
     when "110000011101" => data <= saw_rom(3101);
     when "110000011110" => data <= saw_rom(3102);
     when "110000011111" => data <= saw_rom(3103);
     when "110000100000" => data <= saw_rom(3104);
     when "110000100001" => data <= saw_rom(3105);
     when "110000100010" => data <= saw_rom(3106);
     when "110000100011" => data <= saw_rom(3107);
     when "110000100100" => data <= saw_rom(3108);
     when "110000100101" => data <= saw_rom(3109);
     when "110000100110" => data <= saw_rom(3110);
     when "110000100111" => data <= saw_rom(3111);
     when "110000101000" => data <= saw_rom(3112);
     when "110000101001" => data <= saw_rom(3113);
     when "110000101010" => data <= saw_rom(3114);
     when "110000101011" => data <= saw_rom(3115);
     when "110000101100" => data <= saw_rom(3116);
     when "110000101101" => data <= saw_rom(3117);
     when "110000101110" => data <= saw_rom(3118);
     when "110000101111" => data <= saw_rom(3119);
     when "110000110000" => data <= saw_rom(3120);
     when "110000110001" => data <= saw_rom(3121);
     when "110000110010" => data <= saw_rom(3122);
     when "110000110011" => data <= saw_rom(3123);
     when "110000110100" => data <= saw_rom(3124);
     when "110000110101" => data <= saw_rom(3125);
     when "110000110110" => data <= saw_rom(3126);
     when "110000110111" => data <= saw_rom(3127);
     when "110000111000" => data <= saw_rom(3128);
     when "110000111001" => data <= saw_rom(3129);
     when "110000111010" => data <= saw_rom(3130);
     when "110000111011" => data <= saw_rom(3131);
     when "110000111100" => data <= saw_rom(3132);
     when "110000111101" => data <= saw_rom(3133);
     when "110000111110" => data <= saw_rom(3134);
     when "110000111111" => data <= saw_rom(3135);
     when "110001000000" => data <= saw_rom(3136);
     when "110001000001" => data <= saw_rom(3137);
     when "110001000010" => data <= saw_rom(3138);
     when "110001000011" => data <= saw_rom(3139);
     when "110001000100" => data <= saw_rom(3140);
     when "110001000101" => data <= saw_rom(3141);
     when "110001000110" => data <= saw_rom(3142);
     when "110001000111" => data <= saw_rom(3143);
     when "110001001000" => data <= saw_rom(3144);
     when "110001001001" => data <= saw_rom(3145);
     when "110001001010" => data <= saw_rom(3146);
     when "110001001011" => data <= saw_rom(3147);
     when "110001001100" => data <= saw_rom(3148);
     when "110001001101" => data <= saw_rom(3149);
     when "110001001110" => data <= saw_rom(3150);
     when "110001001111" => data <= saw_rom(3151);
     when "110001010000" => data <= saw_rom(3152);
     when "110001010001" => data <= saw_rom(3153);
     when "110001010010" => data <= saw_rom(3154);
     when "110001010011" => data <= saw_rom(3155);
     when "110001010100" => data <= saw_rom(3156);
     when "110001010101" => data <= saw_rom(3157);
     when "110001010110" => data <= saw_rom(3158);
     when "110001010111" => data <= saw_rom(3159);
     when "110001011000" => data <= saw_rom(3160);
     when "110001011001" => data <= saw_rom(3161);
     when "110001011010" => data <= saw_rom(3162);
     when "110001011011" => data <= saw_rom(3163);
     when "110001011100" => data <= saw_rom(3164);
     when "110001011101" => data <= saw_rom(3165);
     when "110001011110" => data <= saw_rom(3166);
     when "110001011111" => data <= saw_rom(3167);
     when "110001100000" => data <= saw_rom(3168);
     when "110001100001" => data <= saw_rom(3169);
     when "110001100010" => data <= saw_rom(3170);
     when "110001100011" => data <= saw_rom(3171);
     when "110001100100" => data <= saw_rom(3172);
     when "110001100101" => data <= saw_rom(3173);
     when "110001100110" => data <= saw_rom(3174);
     when "110001100111" => data <= saw_rom(3175);
     when "110001101000" => data <= saw_rom(3176);
     when "110001101001" => data <= saw_rom(3177);
     when "110001101010" => data <= saw_rom(3178);
     when "110001101011" => data <= saw_rom(3179);
     when "110001101100" => data <= saw_rom(3180);
     when "110001101101" => data <= saw_rom(3181);
     when "110001101110" => data <= saw_rom(3182);
     when "110001101111" => data <= saw_rom(3183);
     when "110001110000" => data <= saw_rom(3184);
     when "110001110001" => data <= saw_rom(3185);
     when "110001110010" => data <= saw_rom(3186);
     when "110001110011" => data <= saw_rom(3187);
     when "110001110100" => data <= saw_rom(3188);
     when "110001110101" => data <= saw_rom(3189);
     when "110001110110" => data <= saw_rom(3190);
     when "110001110111" => data <= saw_rom(3191);
     when "110001111000" => data <= saw_rom(3192);
     when "110001111001" => data <= saw_rom(3193);
     when "110001111010" => data <= saw_rom(3194);
     when "110001111011" => data <= saw_rom(3195);
     when "110001111100" => data <= saw_rom(3196);
     when "110001111101" => data <= saw_rom(3197);
     when "110001111110" => data <= saw_rom(3198);
     when "110001111111" => data <= saw_rom(3199);
     when "110010000000" => data <= saw_rom(3200);
     when "110010000001" => data <= saw_rom(3201);
     when "110010000010" => data <= saw_rom(3202);
     when "110010000011" => data <= saw_rom(3203);
     when "110010000100" => data <= saw_rom(3204);
     when "110010000101" => data <= saw_rom(3205);
     when "110010000110" => data <= saw_rom(3206);
     when "110010000111" => data <= saw_rom(3207);
     when "110010001000" => data <= saw_rom(3208);
     when "110010001001" => data <= saw_rom(3209);
     when "110010001010" => data <= saw_rom(3210);
     when "110010001011" => data <= saw_rom(3211);
     when "110010001100" => data <= saw_rom(3212);
     when "110010001101" => data <= saw_rom(3213);
     when "110010001110" => data <= saw_rom(3214);
     when "110010001111" => data <= saw_rom(3215);
     when "110010010000" => data <= saw_rom(3216);
     when "110010010001" => data <= saw_rom(3217);
     when "110010010010" => data <= saw_rom(3218);
     when "110010010011" => data <= saw_rom(3219);
     when "110010010100" => data <= saw_rom(3220);
     when "110010010101" => data <= saw_rom(3221);
     when "110010010110" => data <= saw_rom(3222);
     when "110010010111" => data <= saw_rom(3223);
     when "110010011000" => data <= saw_rom(3224);
     when "110010011001" => data <= saw_rom(3225);
     when "110010011010" => data <= saw_rom(3226);
     when "110010011011" => data <= saw_rom(3227);
     when "110010011100" => data <= saw_rom(3228);
     when "110010011101" => data <= saw_rom(3229);
     when "110010011110" => data <= saw_rom(3230);
     when "110010011111" => data <= saw_rom(3231);
     when "110010100000" => data <= saw_rom(3232);
     when "110010100001" => data <= saw_rom(3233);
     when "110010100010" => data <= saw_rom(3234);
     when "110010100011" => data <= saw_rom(3235);
     when "110010100100" => data <= saw_rom(3236);
     when "110010100101" => data <= saw_rom(3237);
     when "110010100110" => data <= saw_rom(3238);
     when "110010100111" => data <= saw_rom(3239);
     when "110010101000" => data <= saw_rom(3240);
     when "110010101001" => data <= saw_rom(3241);
     when "110010101010" => data <= saw_rom(3242);
     when "110010101011" => data <= saw_rom(3243);
     when "110010101100" => data <= saw_rom(3244);
     when "110010101101" => data <= saw_rom(3245);
     when "110010101110" => data <= saw_rom(3246);
     when "110010101111" => data <= saw_rom(3247);
     when "110010110000" => data <= saw_rom(3248);
     when "110010110001" => data <= saw_rom(3249);
     when "110010110010" => data <= saw_rom(3250);
     when "110010110011" => data <= saw_rom(3251);
     when "110010110100" => data <= saw_rom(3252);
     when "110010110101" => data <= saw_rom(3253);
     when "110010110110" => data <= saw_rom(3254);
     when "110010110111" => data <= saw_rom(3255);
     when "110010111000" => data <= saw_rom(3256);
     when "110010111001" => data <= saw_rom(3257);
     when "110010111010" => data <= saw_rom(3258);
     when "110010111011" => data <= saw_rom(3259);
     when "110010111100" => data <= saw_rom(3260);
     when "110010111101" => data <= saw_rom(3261);
     when "110010111110" => data <= saw_rom(3262);
     when "110010111111" => data <= saw_rom(3263);
     when "110011000000" => data <= saw_rom(3264);
     when "110011000001" => data <= saw_rom(3265);
     when "110011000010" => data <= saw_rom(3266);
     when "110011000011" => data <= saw_rom(3267);
     when "110011000100" => data <= saw_rom(3268);
     when "110011000101" => data <= saw_rom(3269);
     when "110011000110" => data <= saw_rom(3270);
     when "110011000111" => data <= saw_rom(3271);
     when "110011001000" => data <= saw_rom(3272);
     when "110011001001" => data <= saw_rom(3273);
     when "110011001010" => data <= saw_rom(3274);
     when "110011001011" => data <= saw_rom(3275);
     when "110011001100" => data <= saw_rom(3276);
     when "110011001101" => data <= saw_rom(3277);
     when "110011001110" => data <= saw_rom(3278);
     when "110011001111" => data <= saw_rom(3279);
     when "110011010000" => data <= saw_rom(3280);
     when "110011010001" => data <= saw_rom(3281);
     when "110011010010" => data <= saw_rom(3282);
     when "110011010011" => data <= saw_rom(3283);
     when "110011010100" => data <= saw_rom(3284);
     when "110011010101" => data <= saw_rom(3285);
     when "110011010110" => data <= saw_rom(3286);
     when "110011010111" => data <= saw_rom(3287);
     when "110011011000" => data <= saw_rom(3288);
     when "110011011001" => data <= saw_rom(3289);
     when "110011011010" => data <= saw_rom(3290);
     when "110011011011" => data <= saw_rom(3291);
     when "110011011100" => data <= saw_rom(3292);
     when "110011011101" => data <= saw_rom(3293);
     when "110011011110" => data <= saw_rom(3294);
     when "110011011111" => data <= saw_rom(3295);
     when "110011100000" => data <= saw_rom(3296);
     when "110011100001" => data <= saw_rom(3297);
     when "110011100010" => data <= saw_rom(3298);
     when "110011100011" => data <= saw_rom(3299);
     when "110011100100" => data <= saw_rom(3300);
     when "110011100101" => data <= saw_rom(3301);
     when "110011100110" => data <= saw_rom(3302);
     when "110011100111" => data <= saw_rom(3303);
     when "110011101000" => data <= saw_rom(3304);
     when "110011101001" => data <= saw_rom(3305);
     when "110011101010" => data <= saw_rom(3306);
     when "110011101011" => data <= saw_rom(3307);
     when "110011101100" => data <= saw_rom(3308);
     when "110011101101" => data <= saw_rom(3309);
     when "110011101110" => data <= saw_rom(3310);
     when "110011101111" => data <= saw_rom(3311);
     when "110011110000" => data <= saw_rom(3312);
     when "110011110001" => data <= saw_rom(3313);
     when "110011110010" => data <= saw_rom(3314);
     when "110011110011" => data <= saw_rom(3315);
     when "110011110100" => data <= saw_rom(3316);
     when "110011110101" => data <= saw_rom(3317);
     when "110011110110" => data <= saw_rom(3318);
     when "110011110111" => data <= saw_rom(3319);
     when "110011111000" => data <= saw_rom(3320);
     when "110011111001" => data <= saw_rom(3321);
     when "110011111010" => data <= saw_rom(3322);
     when "110011111011" => data <= saw_rom(3323);
     when "110011111100" => data <= saw_rom(3324);
     when "110011111101" => data <= saw_rom(3325);
     when "110011111110" => data <= saw_rom(3326);
     when "110011111111" => data <= saw_rom(3327);
     when "110100000000" => data <= saw_rom(3328);
     when "110100000001" => data <= saw_rom(3329);
     when "110100000010" => data <= saw_rom(3330);
     when "110100000011" => data <= saw_rom(3331);
     when "110100000100" => data <= saw_rom(3332);
     when "110100000101" => data <= saw_rom(3333);
     when "110100000110" => data <= saw_rom(3334);
     when "110100000111" => data <= saw_rom(3335);
     when "110100001000" => data <= saw_rom(3336);
     when "110100001001" => data <= saw_rom(3337);
     when "110100001010" => data <= saw_rom(3338);
     when "110100001011" => data <= saw_rom(3339);
     when "110100001100" => data <= saw_rom(3340);
     when "110100001101" => data <= saw_rom(3341);
     when "110100001110" => data <= saw_rom(3342);
     when "110100001111" => data <= saw_rom(3343);
     when "110100010000" => data <= saw_rom(3344);
     when "110100010001" => data <= saw_rom(3345);
     when "110100010010" => data <= saw_rom(3346);
     when "110100010011" => data <= saw_rom(3347);
     when "110100010100" => data <= saw_rom(3348);
     when "110100010101" => data <= saw_rom(3349);
     when "110100010110" => data <= saw_rom(3350);
     when "110100010111" => data <= saw_rom(3351);
     when "110100011000" => data <= saw_rom(3352);
     when "110100011001" => data <= saw_rom(3353);
     when "110100011010" => data <= saw_rom(3354);
     when "110100011011" => data <= saw_rom(3355);
     when "110100011100" => data <= saw_rom(3356);
     when "110100011101" => data <= saw_rom(3357);
     when "110100011110" => data <= saw_rom(3358);
     when "110100011111" => data <= saw_rom(3359);
     when "110100100000" => data <= saw_rom(3360);
     when "110100100001" => data <= saw_rom(3361);
     when "110100100010" => data <= saw_rom(3362);
     when "110100100011" => data <= saw_rom(3363);
     when "110100100100" => data <= saw_rom(3364);
     when "110100100101" => data <= saw_rom(3365);
     when "110100100110" => data <= saw_rom(3366);
     when "110100100111" => data <= saw_rom(3367);
     when "110100101000" => data <= saw_rom(3368);
     when "110100101001" => data <= saw_rom(3369);
     when "110100101010" => data <= saw_rom(3370);
     when "110100101011" => data <= saw_rom(3371);
     when "110100101100" => data <= saw_rom(3372);
     when "110100101101" => data <= saw_rom(3373);
     when "110100101110" => data <= saw_rom(3374);
     when "110100101111" => data <= saw_rom(3375);
     when "110100110000" => data <= saw_rom(3376);
     when "110100110001" => data <= saw_rom(3377);
     when "110100110010" => data <= saw_rom(3378);
     when "110100110011" => data <= saw_rom(3379);
     when "110100110100" => data <= saw_rom(3380);
     when "110100110101" => data <= saw_rom(3381);
     when "110100110110" => data <= saw_rom(3382);
     when "110100110111" => data <= saw_rom(3383);
     when "110100111000" => data <= saw_rom(3384);
     when "110100111001" => data <= saw_rom(3385);
     when "110100111010" => data <= saw_rom(3386);
     when "110100111011" => data <= saw_rom(3387);
     when "110100111100" => data <= saw_rom(3388);
     when "110100111101" => data <= saw_rom(3389);
     when "110100111110" => data <= saw_rom(3390);
     when "110100111111" => data <= saw_rom(3391);
     when "110101000000" => data <= saw_rom(3392);
     when "110101000001" => data <= saw_rom(3393);
     when "110101000010" => data <= saw_rom(3394);
     when "110101000011" => data <= saw_rom(3395);
     when "110101000100" => data <= saw_rom(3396);
     when "110101000101" => data <= saw_rom(3397);
     when "110101000110" => data <= saw_rom(3398);
     when "110101000111" => data <= saw_rom(3399);
     when "110101001000" => data <= saw_rom(3400);
     when "110101001001" => data <= saw_rom(3401);
     when "110101001010" => data <= saw_rom(3402);
     when "110101001011" => data <= saw_rom(3403);
     when "110101001100" => data <= saw_rom(3404);
     when "110101001101" => data <= saw_rom(3405);
     when "110101001110" => data <= saw_rom(3406);
     when "110101001111" => data <= saw_rom(3407);
     when "110101010000" => data <= saw_rom(3408);
     when "110101010001" => data <= saw_rom(3409);
     when "110101010010" => data <= saw_rom(3410);
     when "110101010011" => data <= saw_rom(3411);
     when "110101010100" => data <= saw_rom(3412);
     when "110101010101" => data <= saw_rom(3413);
     when "110101010110" => data <= saw_rom(3414);
     when "110101010111" => data <= saw_rom(3415);
     when "110101011000" => data <= saw_rom(3416);
     when "110101011001" => data <= saw_rom(3417);
     when "110101011010" => data <= saw_rom(3418);
     when "110101011011" => data <= saw_rom(3419);
     when "110101011100" => data <= saw_rom(3420);
     when "110101011101" => data <= saw_rom(3421);
     when "110101011110" => data <= saw_rom(3422);
     when "110101011111" => data <= saw_rom(3423);
     when "110101100000" => data <= saw_rom(3424);
     when "110101100001" => data <= saw_rom(3425);
     when "110101100010" => data <= saw_rom(3426);
     when "110101100011" => data <= saw_rom(3427);
     when "110101100100" => data <= saw_rom(3428);
     when "110101100101" => data <= saw_rom(3429);
     when "110101100110" => data <= saw_rom(3430);
     when "110101100111" => data <= saw_rom(3431);
     when "110101101000" => data <= saw_rom(3432);
     when "110101101001" => data <= saw_rom(3433);
     when "110101101010" => data <= saw_rom(3434);
     when "110101101011" => data <= saw_rom(3435);
     when "110101101100" => data <= saw_rom(3436);
     when "110101101101" => data <= saw_rom(3437);
     when "110101101110" => data <= saw_rom(3438);
     when "110101101111" => data <= saw_rom(3439);
     when "110101110000" => data <= saw_rom(3440);
     when "110101110001" => data <= saw_rom(3441);
     when "110101110010" => data <= saw_rom(3442);
     when "110101110011" => data <= saw_rom(3443);
     when "110101110100" => data <= saw_rom(3444);
     when "110101110101" => data <= saw_rom(3445);
     when "110101110110" => data <= saw_rom(3446);
     when "110101110111" => data <= saw_rom(3447);
     when "110101111000" => data <= saw_rom(3448);
     when "110101111001" => data <= saw_rom(3449);
     when "110101111010" => data <= saw_rom(3450);
     when "110101111011" => data <= saw_rom(3451);
     when "110101111100" => data <= saw_rom(3452);
     when "110101111101" => data <= saw_rom(3453);
     when "110101111110" => data <= saw_rom(3454);
     when "110101111111" => data <= saw_rom(3455);
     when "110110000000" => data <= saw_rom(3456);
     when "110110000001" => data <= saw_rom(3457);
     when "110110000010" => data <= saw_rom(3458);
     when "110110000011" => data <= saw_rom(3459);
     when "110110000100" => data <= saw_rom(3460);
     when "110110000101" => data <= saw_rom(3461);
     when "110110000110" => data <= saw_rom(3462);
     when "110110000111" => data <= saw_rom(3463);
     when "110110001000" => data <= saw_rom(3464);
     when "110110001001" => data <= saw_rom(3465);
     when "110110001010" => data <= saw_rom(3466);
     when "110110001011" => data <= saw_rom(3467);
     when "110110001100" => data <= saw_rom(3468);
     when "110110001101" => data <= saw_rom(3469);
     when "110110001110" => data <= saw_rom(3470);
     when "110110001111" => data <= saw_rom(3471);
     when "110110010000" => data <= saw_rom(3472);
     when "110110010001" => data <= saw_rom(3473);
     when "110110010010" => data <= saw_rom(3474);
     when "110110010011" => data <= saw_rom(3475);
     when "110110010100" => data <= saw_rom(3476);
     when "110110010101" => data <= saw_rom(3477);
     when "110110010110" => data <= saw_rom(3478);
     when "110110010111" => data <= saw_rom(3479);
     when "110110011000" => data <= saw_rom(3480);
     when "110110011001" => data <= saw_rom(3481);
     when "110110011010" => data <= saw_rom(3482);
     when "110110011011" => data <= saw_rom(3483);
     when "110110011100" => data <= saw_rom(3484);
     when "110110011101" => data <= saw_rom(3485);
     when "110110011110" => data <= saw_rom(3486);
     when "110110011111" => data <= saw_rom(3487);
     when "110110100000" => data <= saw_rom(3488);
     when "110110100001" => data <= saw_rom(3489);
     when "110110100010" => data <= saw_rom(3490);
     when "110110100011" => data <= saw_rom(3491);
     when "110110100100" => data <= saw_rom(3492);
     when "110110100101" => data <= saw_rom(3493);
     when "110110100110" => data <= saw_rom(3494);
     when "110110100111" => data <= saw_rom(3495);
     when "110110101000" => data <= saw_rom(3496);
     when "110110101001" => data <= saw_rom(3497);
     when "110110101010" => data <= saw_rom(3498);
     when "110110101011" => data <= saw_rom(3499);
     when "110110101100" => data <= saw_rom(3500);
     when "110110101101" => data <= saw_rom(3501);
     when "110110101110" => data <= saw_rom(3502);
     when "110110101111" => data <= saw_rom(3503);
     when "110110110000" => data <= saw_rom(3504);
     when "110110110001" => data <= saw_rom(3505);
     when "110110110010" => data <= saw_rom(3506);
     when "110110110011" => data <= saw_rom(3507);
     when "110110110100" => data <= saw_rom(3508);
     when "110110110101" => data <= saw_rom(3509);
     when "110110110110" => data <= saw_rom(3510);
     when "110110110111" => data <= saw_rom(3511);
     when "110110111000" => data <= saw_rom(3512);
     when "110110111001" => data <= saw_rom(3513);
     when "110110111010" => data <= saw_rom(3514);
     when "110110111011" => data <= saw_rom(3515);
     when "110110111100" => data <= saw_rom(3516);
     when "110110111101" => data <= saw_rom(3517);
     when "110110111110" => data <= saw_rom(3518);
     when "110110111111" => data <= saw_rom(3519);
     when "110111000000" => data <= saw_rom(3520);
     when "110111000001" => data <= saw_rom(3521);
     when "110111000010" => data <= saw_rom(3522);
     when "110111000011" => data <= saw_rom(3523);
     when "110111000100" => data <= saw_rom(3524);
     when "110111000101" => data <= saw_rom(3525);
     when "110111000110" => data <= saw_rom(3526);
     when "110111000111" => data <= saw_rom(3527);
     when "110111001000" => data <= saw_rom(3528);
     when "110111001001" => data <= saw_rom(3529);
     when "110111001010" => data <= saw_rom(3530);
     when "110111001011" => data <= saw_rom(3531);
     when "110111001100" => data <= saw_rom(3532);
     when "110111001101" => data <= saw_rom(3533);
     when "110111001110" => data <= saw_rom(3534);
     when "110111001111" => data <= saw_rom(3535);
     when "110111010000" => data <= saw_rom(3536);
     when "110111010001" => data <= saw_rom(3537);
     when "110111010010" => data <= saw_rom(3538);
     when "110111010011" => data <= saw_rom(3539);
     when "110111010100" => data <= saw_rom(3540);
     when "110111010101" => data <= saw_rom(3541);
     when "110111010110" => data <= saw_rom(3542);
     when "110111010111" => data <= saw_rom(3543);
     when "110111011000" => data <= saw_rom(3544);
     when "110111011001" => data <= saw_rom(3545);
     when "110111011010" => data <= saw_rom(3546);
     when "110111011011" => data <= saw_rom(3547);
     when "110111011100" => data <= saw_rom(3548);
     when "110111011101" => data <= saw_rom(3549);
     when "110111011110" => data <= saw_rom(3550);
     when "110111011111" => data <= saw_rom(3551);
     when "110111100000" => data <= saw_rom(3552);
     when "110111100001" => data <= saw_rom(3553);
     when "110111100010" => data <= saw_rom(3554);
     when "110111100011" => data <= saw_rom(3555);
     when "110111100100" => data <= saw_rom(3556);
     when "110111100101" => data <= saw_rom(3557);
     when "110111100110" => data <= saw_rom(3558);
     when "110111100111" => data <= saw_rom(3559);
     when "110111101000" => data <= saw_rom(3560);
     when "110111101001" => data <= saw_rom(3561);
     when "110111101010" => data <= saw_rom(3562);
     when "110111101011" => data <= saw_rom(3563);
     when "110111101100" => data <= saw_rom(3564);
     when "110111101101" => data <= saw_rom(3565);
     when "110111101110" => data <= saw_rom(3566);
     when "110111101111" => data <= saw_rom(3567);
     when "110111110000" => data <= saw_rom(3568);
     when "110111110001" => data <= saw_rom(3569);
     when "110111110010" => data <= saw_rom(3570);
     when "110111110011" => data <= saw_rom(3571);
     when "110111110100" => data <= saw_rom(3572);
     when "110111110101" => data <= saw_rom(3573);
     when "110111110110" => data <= saw_rom(3574);
     when "110111110111" => data <= saw_rom(3575);
     when "110111111000" => data <= saw_rom(3576);
     when "110111111001" => data <= saw_rom(3577);
     when "110111111010" => data <= saw_rom(3578);
     when "110111111011" => data <= saw_rom(3579);
     when "110111111100" => data <= saw_rom(3580);
     when "110111111101" => data <= saw_rom(3581);
     when "110111111110" => data <= saw_rom(3582);
     when "110111111111" => data <= saw_rom(3583);
     when "111000000000" => data <= saw_rom(3584);
     when "111000000001" => data <= saw_rom(3585);
     when "111000000010" => data <= saw_rom(3586);
     when "111000000011" => data <= saw_rom(3587);
     when "111000000100" => data <= saw_rom(3588);
     when "111000000101" => data <= saw_rom(3589);
     when "111000000110" => data <= saw_rom(3590);
     when "111000000111" => data <= saw_rom(3591);
     when "111000001000" => data <= saw_rom(3592);
     when "111000001001" => data <= saw_rom(3593);
     when "111000001010" => data <= saw_rom(3594);
     when "111000001011" => data <= saw_rom(3595);
     when "111000001100" => data <= saw_rom(3596);
     when "111000001101" => data <= saw_rom(3597);
     when "111000001110" => data <= saw_rom(3598);
     when "111000001111" => data <= saw_rom(3599);
     when "111000010000" => data <= saw_rom(3600);
     when "111000010001" => data <= saw_rom(3601);
     when "111000010010" => data <= saw_rom(3602);
     when "111000010011" => data <= saw_rom(3603);
     when "111000010100" => data <= saw_rom(3604);
     when "111000010101" => data <= saw_rom(3605);
     when "111000010110" => data <= saw_rom(3606);
     when "111000010111" => data <= saw_rom(3607);
     when "111000011000" => data <= saw_rom(3608);
     when "111000011001" => data <= saw_rom(3609);
     when "111000011010" => data <= saw_rom(3610);
     when "111000011011" => data <= saw_rom(3611);
     when "111000011100" => data <= saw_rom(3612);
     when "111000011101" => data <= saw_rom(3613);
     when "111000011110" => data <= saw_rom(3614);
     when "111000011111" => data <= saw_rom(3615);
     when "111000100000" => data <= saw_rom(3616);
     when "111000100001" => data <= saw_rom(3617);
     when "111000100010" => data <= saw_rom(3618);
     when "111000100011" => data <= saw_rom(3619);
     when "111000100100" => data <= saw_rom(3620);
     when "111000100101" => data <= saw_rom(3621);
     when "111000100110" => data <= saw_rom(3622);
     when "111000100111" => data <= saw_rom(3623);
     when "111000101000" => data <= saw_rom(3624);
     when "111000101001" => data <= saw_rom(3625);
     when "111000101010" => data <= saw_rom(3626);
     when "111000101011" => data <= saw_rom(3627);
     when "111000101100" => data <= saw_rom(3628);
     when "111000101101" => data <= saw_rom(3629);
     when "111000101110" => data <= saw_rom(3630);
     when "111000101111" => data <= saw_rom(3631);
     when "111000110000" => data <= saw_rom(3632);
     when "111000110001" => data <= saw_rom(3633);
     when "111000110010" => data <= saw_rom(3634);
     when "111000110011" => data <= saw_rom(3635);
     when "111000110100" => data <= saw_rom(3636);
     when "111000110101" => data <= saw_rom(3637);
     when "111000110110" => data <= saw_rom(3638);
     when "111000110111" => data <= saw_rom(3639);
     when "111000111000" => data <= saw_rom(3640);
     when "111000111001" => data <= saw_rom(3641);
     when "111000111010" => data <= saw_rom(3642);
     when "111000111011" => data <= saw_rom(3643);
     when "111000111100" => data <= saw_rom(3644);
     when "111000111101" => data <= saw_rom(3645);
     when "111000111110" => data <= saw_rom(3646);
     when "111000111111" => data <= saw_rom(3647);
     when "111001000000" => data <= saw_rom(3648);
     when "111001000001" => data <= saw_rom(3649);
     when "111001000010" => data <= saw_rom(3650);
     when "111001000011" => data <= saw_rom(3651);
     when "111001000100" => data <= saw_rom(3652);
     when "111001000101" => data <= saw_rom(3653);
     when "111001000110" => data <= saw_rom(3654);
     when "111001000111" => data <= saw_rom(3655);
     when "111001001000" => data <= saw_rom(3656);
     when "111001001001" => data <= saw_rom(3657);
     when "111001001010" => data <= saw_rom(3658);
     when "111001001011" => data <= saw_rom(3659);
     when "111001001100" => data <= saw_rom(3660);
     when "111001001101" => data <= saw_rom(3661);
     when "111001001110" => data <= saw_rom(3662);
     when "111001001111" => data <= saw_rom(3663);
     when "111001010000" => data <= saw_rom(3664);
     when "111001010001" => data <= saw_rom(3665);
     when "111001010010" => data <= saw_rom(3666);
     when "111001010011" => data <= saw_rom(3667);
     when "111001010100" => data <= saw_rom(3668);
     when "111001010101" => data <= saw_rom(3669);
     when "111001010110" => data <= saw_rom(3670);
     when "111001010111" => data <= saw_rom(3671);
     when "111001011000" => data <= saw_rom(3672);
     when "111001011001" => data <= saw_rom(3673);
     when "111001011010" => data <= saw_rom(3674);
     when "111001011011" => data <= saw_rom(3675);
     when "111001011100" => data <= saw_rom(3676);
     when "111001011101" => data <= saw_rom(3677);
     when "111001011110" => data <= saw_rom(3678);
     when "111001011111" => data <= saw_rom(3679);
     when "111001100000" => data <= saw_rom(3680);
     when "111001100001" => data <= saw_rom(3681);
     when "111001100010" => data <= saw_rom(3682);
     when "111001100011" => data <= saw_rom(3683);
     when "111001100100" => data <= saw_rom(3684);
     when "111001100101" => data <= saw_rom(3685);
     when "111001100110" => data <= saw_rom(3686);
     when "111001100111" => data <= saw_rom(3687);
     when "111001101000" => data <= saw_rom(3688);
     when "111001101001" => data <= saw_rom(3689);
     when "111001101010" => data <= saw_rom(3690);
     when "111001101011" => data <= saw_rom(3691);
     when "111001101100" => data <= saw_rom(3692);
     when "111001101101" => data <= saw_rom(3693);
     when "111001101110" => data <= saw_rom(3694);
     when "111001101111" => data <= saw_rom(3695);
     when "111001110000" => data <= saw_rom(3696);
     when "111001110001" => data <= saw_rom(3697);
     when "111001110010" => data <= saw_rom(3698);
     when "111001110011" => data <= saw_rom(3699);
     when "111001110100" => data <= saw_rom(3700);
     when "111001110101" => data <= saw_rom(3701);
     when "111001110110" => data <= saw_rom(3702);
     when "111001110111" => data <= saw_rom(3703);
     when "111001111000" => data <= saw_rom(3704);
     when "111001111001" => data <= saw_rom(3705);
     when "111001111010" => data <= saw_rom(3706);
     when "111001111011" => data <= saw_rom(3707);
     when "111001111100" => data <= saw_rom(3708);
     when "111001111101" => data <= saw_rom(3709);
     when "111001111110" => data <= saw_rom(3710);
     when "111001111111" => data <= saw_rom(3711);
     when "111010000000" => data <= saw_rom(3712);
     when "111010000001" => data <= saw_rom(3713);
     when "111010000010" => data <= saw_rom(3714);
     when "111010000011" => data <= saw_rom(3715);
     when "111010000100" => data <= saw_rom(3716);
     when "111010000101" => data <= saw_rom(3717);
     when "111010000110" => data <= saw_rom(3718);
     when "111010000111" => data <= saw_rom(3719);
     when "111010001000" => data <= saw_rom(3720);
     when "111010001001" => data <= saw_rom(3721);
     when "111010001010" => data <= saw_rom(3722);
     when "111010001011" => data <= saw_rom(3723);
     when "111010001100" => data <= saw_rom(3724);
     when "111010001101" => data <= saw_rom(3725);
     when "111010001110" => data <= saw_rom(3726);
     when "111010001111" => data <= saw_rom(3727);
     when "111010010000" => data <= saw_rom(3728);
     when "111010010001" => data <= saw_rom(3729);
     when "111010010010" => data <= saw_rom(3730);
     when "111010010011" => data <= saw_rom(3731);
     when "111010010100" => data <= saw_rom(3732);
     when "111010010101" => data <= saw_rom(3733);
     when "111010010110" => data <= saw_rom(3734);
     when "111010010111" => data <= saw_rom(3735);
     when "111010011000" => data <= saw_rom(3736);
     when "111010011001" => data <= saw_rom(3737);
     when "111010011010" => data <= saw_rom(3738);
     when "111010011011" => data <= saw_rom(3739);
     when "111010011100" => data <= saw_rom(3740);
     when "111010011101" => data <= saw_rom(3741);
     when "111010011110" => data <= saw_rom(3742);
     when "111010011111" => data <= saw_rom(3743);
     when "111010100000" => data <= saw_rom(3744);
     when "111010100001" => data <= saw_rom(3745);
     when "111010100010" => data <= saw_rom(3746);
     when "111010100011" => data <= saw_rom(3747);
     when "111010100100" => data <= saw_rom(3748);
     when "111010100101" => data <= saw_rom(3749);
     when "111010100110" => data <= saw_rom(3750);
     when "111010100111" => data <= saw_rom(3751);
     when "111010101000" => data <= saw_rom(3752);
     when "111010101001" => data <= saw_rom(3753);
     when "111010101010" => data <= saw_rom(3754);
     when "111010101011" => data <= saw_rom(3755);
     when "111010101100" => data <= saw_rom(3756);
     when "111010101101" => data <= saw_rom(3757);
     when "111010101110" => data <= saw_rom(3758);
     when "111010101111" => data <= saw_rom(3759);
     when "111010110000" => data <= saw_rom(3760);
     when "111010110001" => data <= saw_rom(3761);
     when "111010110010" => data <= saw_rom(3762);
     when "111010110011" => data <= saw_rom(3763);
     when "111010110100" => data <= saw_rom(3764);
     when "111010110101" => data <= saw_rom(3765);
     when "111010110110" => data <= saw_rom(3766);
     when "111010110111" => data <= saw_rom(3767);
     when "111010111000" => data <= saw_rom(3768);
     when "111010111001" => data <= saw_rom(3769);
     when "111010111010" => data <= saw_rom(3770);
     when "111010111011" => data <= saw_rom(3771);
     when "111010111100" => data <= saw_rom(3772);
     when "111010111101" => data <= saw_rom(3773);
     when "111010111110" => data <= saw_rom(3774);
     when "111010111111" => data <= saw_rom(3775);
     when "111011000000" => data <= saw_rom(3776);
     when "111011000001" => data <= saw_rom(3777);
     when "111011000010" => data <= saw_rom(3778);
     when "111011000011" => data <= saw_rom(3779);
     when "111011000100" => data <= saw_rom(3780);
     when "111011000101" => data <= saw_rom(3781);
     when "111011000110" => data <= saw_rom(3782);
     when "111011000111" => data <= saw_rom(3783);
     when "111011001000" => data <= saw_rom(3784);
     when "111011001001" => data <= saw_rom(3785);
     when "111011001010" => data <= saw_rom(3786);
     when "111011001011" => data <= saw_rom(3787);
     when "111011001100" => data <= saw_rom(3788);
     when "111011001101" => data <= saw_rom(3789);
     when "111011001110" => data <= saw_rom(3790);
     when "111011001111" => data <= saw_rom(3791);
     when "111011010000" => data <= saw_rom(3792);
     when "111011010001" => data <= saw_rom(3793);
     when "111011010010" => data <= saw_rom(3794);
     when "111011010011" => data <= saw_rom(3795);
     when "111011010100" => data <= saw_rom(3796);
     when "111011010101" => data <= saw_rom(3797);
     when "111011010110" => data <= saw_rom(3798);
     when "111011010111" => data <= saw_rom(3799);
     when "111011011000" => data <= saw_rom(3800);
     when "111011011001" => data <= saw_rom(3801);
     when "111011011010" => data <= saw_rom(3802);
     when "111011011011" => data <= saw_rom(3803);
     when "111011011100" => data <= saw_rom(3804);
     when "111011011101" => data <= saw_rom(3805);
     when "111011011110" => data <= saw_rom(3806);
     when "111011011111" => data <= saw_rom(3807);
     when "111011100000" => data <= saw_rom(3808);
     when "111011100001" => data <= saw_rom(3809);
     when "111011100010" => data <= saw_rom(3810);
     when "111011100011" => data <= saw_rom(3811);
     when "111011100100" => data <= saw_rom(3812);
     when "111011100101" => data <= saw_rom(3813);
     when "111011100110" => data <= saw_rom(3814);
     when "111011100111" => data <= saw_rom(3815);
     when "111011101000" => data <= saw_rom(3816);
     when "111011101001" => data <= saw_rom(3817);
     when "111011101010" => data <= saw_rom(3818);
     when "111011101011" => data <= saw_rom(3819);
     when "111011101100" => data <= saw_rom(3820);
     when "111011101101" => data <= saw_rom(3821);
     when "111011101110" => data <= saw_rom(3822);
     when "111011101111" => data <= saw_rom(3823);
     when "111011110000" => data <= saw_rom(3824);
     when "111011110001" => data <= saw_rom(3825);
     when "111011110010" => data <= saw_rom(3826);
     when "111011110011" => data <= saw_rom(3827);
     when "111011110100" => data <= saw_rom(3828);
     when "111011110101" => data <= saw_rom(3829);
     when "111011110110" => data <= saw_rom(3830);
     when "111011110111" => data <= saw_rom(3831);
     when "111011111000" => data <= saw_rom(3832);
     when "111011111001" => data <= saw_rom(3833);
     when "111011111010" => data <= saw_rom(3834);
     when "111011111011" => data <= saw_rom(3835);
     when "111011111100" => data <= saw_rom(3836);
     when "111011111101" => data <= saw_rom(3837);
     when "111011111110" => data <= saw_rom(3838);
     when "111011111111" => data <= saw_rom(3839);
     when "111100000000" => data <= saw_rom(3840);
     when "111100000001" => data <= saw_rom(3841);
     when "111100000010" => data <= saw_rom(3842);
     when "111100000011" => data <= saw_rom(3843);
     when "111100000100" => data <= saw_rom(3844);
     when "111100000101" => data <= saw_rom(3845);
     when "111100000110" => data <= saw_rom(3846);
     when "111100000111" => data <= saw_rom(3847);
     when "111100001000" => data <= saw_rom(3848);
     when "111100001001" => data <= saw_rom(3849);
     when "111100001010" => data <= saw_rom(3850);
     when "111100001011" => data <= saw_rom(3851);
     when "111100001100" => data <= saw_rom(3852);
     when "111100001101" => data <= saw_rom(3853);
     when "111100001110" => data <= saw_rom(3854);
     when "111100001111" => data <= saw_rom(3855);
     when "111100010000" => data <= saw_rom(3856);
     when "111100010001" => data <= saw_rom(3857);
     when "111100010010" => data <= saw_rom(3858);
     when "111100010011" => data <= saw_rom(3859);
     when "111100010100" => data <= saw_rom(3860);
     when "111100010101" => data <= saw_rom(3861);
     when "111100010110" => data <= saw_rom(3862);
     when "111100010111" => data <= saw_rom(3863);
     when "111100011000" => data <= saw_rom(3864);
     when "111100011001" => data <= saw_rom(3865);
     when "111100011010" => data <= saw_rom(3866);
     when "111100011011" => data <= saw_rom(3867);
     when "111100011100" => data <= saw_rom(3868);
     when "111100011101" => data <= saw_rom(3869);
     when "111100011110" => data <= saw_rom(3870);
     when "111100011111" => data <= saw_rom(3871);
     when "111100100000" => data <= saw_rom(3872);
     when "111100100001" => data <= saw_rom(3873);
     when "111100100010" => data <= saw_rom(3874);
     when "111100100011" => data <= saw_rom(3875);
     when "111100100100" => data <= saw_rom(3876);
     when "111100100101" => data <= saw_rom(3877);
     when "111100100110" => data <= saw_rom(3878);
     when "111100100111" => data <= saw_rom(3879);
     when "111100101000" => data <= saw_rom(3880);
     when "111100101001" => data <= saw_rom(3881);
     when "111100101010" => data <= saw_rom(3882);
     when "111100101011" => data <= saw_rom(3883);
     when "111100101100" => data <= saw_rom(3884);
     when "111100101101" => data <= saw_rom(3885);
     when "111100101110" => data <= saw_rom(3886);
     when "111100101111" => data <= saw_rom(3887);
     when "111100110000" => data <= saw_rom(3888);
     when "111100110001" => data <= saw_rom(3889);
     when "111100110010" => data <= saw_rom(3890);
     when "111100110011" => data <= saw_rom(3891);
     when "111100110100" => data <= saw_rom(3892);
     when "111100110101" => data <= saw_rom(3893);
     when "111100110110" => data <= saw_rom(3894);
     when "111100110111" => data <= saw_rom(3895);
     when "111100111000" => data <= saw_rom(3896);
     when "111100111001" => data <= saw_rom(3897);
     when "111100111010" => data <= saw_rom(3898);
     when "111100111011" => data <= saw_rom(3899);
     when "111100111100" => data <= saw_rom(3900);
     when "111100111101" => data <= saw_rom(3901);
     when "111100111110" => data <= saw_rom(3902);
     when "111100111111" => data <= saw_rom(3903);
     when "111101000000" => data <= saw_rom(3904);
     when "111101000001" => data <= saw_rom(3905);
     when "111101000010" => data <= saw_rom(3906);
     when "111101000011" => data <= saw_rom(3907);
     when "111101000100" => data <= saw_rom(3908);
     when "111101000101" => data <= saw_rom(3909);
     when "111101000110" => data <= saw_rom(3910);
     when "111101000111" => data <= saw_rom(3911);
     when "111101001000" => data <= saw_rom(3912);
     when "111101001001" => data <= saw_rom(3913);
     when "111101001010" => data <= saw_rom(3914);
     when "111101001011" => data <= saw_rom(3915);
     when "111101001100" => data <= saw_rom(3916);
     when "111101001101" => data <= saw_rom(3917);
     when "111101001110" => data <= saw_rom(3918);
     when "111101001111" => data <= saw_rom(3919);
     when "111101010000" => data <= saw_rom(3920);
     when "111101010001" => data <= saw_rom(3921);
     when "111101010010" => data <= saw_rom(3922);
     when "111101010011" => data <= saw_rom(3923);
     when "111101010100" => data <= saw_rom(3924);
     when "111101010101" => data <= saw_rom(3925);
     when "111101010110" => data <= saw_rom(3926);
     when "111101010111" => data <= saw_rom(3927);
     when "111101011000" => data <= saw_rom(3928);
     when "111101011001" => data <= saw_rom(3929);
     when "111101011010" => data <= saw_rom(3930);
     when "111101011011" => data <= saw_rom(3931);
     when "111101011100" => data <= saw_rom(3932);
     when "111101011101" => data <= saw_rom(3933);
     when "111101011110" => data <= saw_rom(3934);
     when "111101011111" => data <= saw_rom(3935);
     when "111101100000" => data <= saw_rom(3936);
     when "111101100001" => data <= saw_rom(3937);
     when "111101100010" => data <= saw_rom(3938);
     when "111101100011" => data <= saw_rom(3939);
     when "111101100100" => data <= saw_rom(3940);
     when "111101100101" => data <= saw_rom(3941);
     when "111101100110" => data <= saw_rom(3942);
     when "111101100111" => data <= saw_rom(3943);
     when "111101101000" => data <= saw_rom(3944);
     when "111101101001" => data <= saw_rom(3945);
     when "111101101010" => data <= saw_rom(3946);
     when "111101101011" => data <= saw_rom(3947);
     when "111101101100" => data <= saw_rom(3948);
     when "111101101101" => data <= saw_rom(3949);
     when "111101101110" => data <= saw_rom(3950);
     when "111101101111" => data <= saw_rom(3951);
     when "111101110000" => data <= saw_rom(3952);
     when "111101110001" => data <= saw_rom(3953);
     when "111101110010" => data <= saw_rom(3954);
     when "111101110011" => data <= saw_rom(3955);
     when "111101110100" => data <= saw_rom(3956);
     when "111101110101" => data <= saw_rom(3957);
     when "111101110110" => data <= saw_rom(3958);
     when "111101110111" => data <= saw_rom(3959);
     when "111101111000" => data <= saw_rom(3960);
     when "111101111001" => data <= saw_rom(3961);
     when "111101111010" => data <= saw_rom(3962);
     when "111101111011" => data <= saw_rom(3963);
     when "111101111100" => data <= saw_rom(3964);
     when "111101111101" => data <= saw_rom(3965);
     when "111101111110" => data <= saw_rom(3966);
     when "111101111111" => data <= saw_rom(3967);
     when "111110000000" => data <= saw_rom(3968);
     when "111110000001" => data <= saw_rom(3969);
     when "111110000010" => data <= saw_rom(3970);
     when "111110000011" => data <= saw_rom(3971);
     when "111110000100" => data <= saw_rom(3972);
     when "111110000101" => data <= saw_rom(3973);
     when "111110000110" => data <= saw_rom(3974);
     when "111110000111" => data <= saw_rom(3975);
     when "111110001000" => data <= saw_rom(3976);
     when "111110001001" => data <= saw_rom(3977);
     when "111110001010" => data <= saw_rom(3978);
     when "111110001011" => data <= saw_rom(3979);
     when "111110001100" => data <= saw_rom(3980);
     when "111110001101" => data <= saw_rom(3981);
     when "111110001110" => data <= saw_rom(3982);
     when "111110001111" => data <= saw_rom(3983);
     when "111110010000" => data <= saw_rom(3984);
     when "111110010001" => data <= saw_rom(3985);
     when "111110010010" => data <= saw_rom(3986);
     when "111110010011" => data <= saw_rom(3987);
     when "111110010100" => data <= saw_rom(3988);
     when "111110010101" => data <= saw_rom(3989);
     when "111110010110" => data <= saw_rom(3990);
     when "111110010111" => data <= saw_rom(3991);
     when "111110011000" => data <= saw_rom(3992);
     when "111110011001" => data <= saw_rom(3993);
     when "111110011010" => data <= saw_rom(3994);
     when "111110011011" => data <= saw_rom(3995);
     when "111110011100" => data <= saw_rom(3996);
     when "111110011101" => data <= saw_rom(3997);
     when "111110011110" => data <= saw_rom(3998);
     when "111110011111" => data <= saw_rom(3999);
     when "111110100000" => data <= saw_rom(4000);
     when "111110100001" => data <= saw_rom(4001);
     when "111110100010" => data <= saw_rom(4002);
     when "111110100011" => data <= saw_rom(4003);
     when "111110100100" => data <= saw_rom(4004);
     when "111110100101" => data <= saw_rom(4005);
     when "111110100110" => data <= saw_rom(4006);
     when "111110100111" => data <= saw_rom(4007);
     when "111110101000" => data <= saw_rom(4008);
     when "111110101001" => data <= saw_rom(4009);
     when "111110101010" => data <= saw_rom(4010);
     when "111110101011" => data <= saw_rom(4011);
     when "111110101100" => data <= saw_rom(4012);
     when "111110101101" => data <= saw_rom(4013);
     when "111110101110" => data <= saw_rom(4014);
     when "111110101111" => data <= saw_rom(4015);
     when "111110110000" => data <= saw_rom(4016);
     when "111110110001" => data <= saw_rom(4017);
     when "111110110010" => data <= saw_rom(4018);
     when "111110110011" => data <= saw_rom(4019);
     when "111110110100" => data <= saw_rom(4020);
     when "111110110101" => data <= saw_rom(4021);
     when "111110110110" => data <= saw_rom(4022);
     when "111110110111" => data <= saw_rom(4023);
     when "111110111000" => data <= saw_rom(4024);
     when "111110111001" => data <= saw_rom(4025);
     when "111110111010" => data <= saw_rom(4026);
     when "111110111011" => data <= saw_rom(4027);
     when "111110111100" => data <= saw_rom(4028);
     when "111110111101" => data <= saw_rom(4029);
     when "111110111110" => data <= saw_rom(4030);
     when "111110111111" => data <= saw_rom(4031);
     when "111111000000" => data <= saw_rom(4032);
     when "111111000001" => data <= saw_rom(4033);
     when "111111000010" => data <= saw_rom(4034);
     when "111111000011" => data <= saw_rom(4035);
     when "111111000100" => data <= saw_rom(4036);
     when "111111000101" => data <= saw_rom(4037);
     when "111111000110" => data <= saw_rom(4038);
     when "111111000111" => data <= saw_rom(4039);
     when "111111001000" => data <= saw_rom(4040);
     when "111111001001" => data <= saw_rom(4041);
     when "111111001010" => data <= saw_rom(4042);
     when "111111001011" => data <= saw_rom(4043);
     when "111111001100" => data <= saw_rom(4044);
     when "111111001101" => data <= saw_rom(4045);
     when "111111001110" => data <= saw_rom(4046);
     when "111111001111" => data <= saw_rom(4047);
     when "111111010000" => data <= saw_rom(4048);
     when "111111010001" => data <= saw_rom(4049);
     when "111111010010" => data <= saw_rom(4050);
     when "111111010011" => data <= saw_rom(4051);
     when "111111010100" => data <= saw_rom(4052);
     when "111111010101" => data <= saw_rom(4053);
     when "111111010110" => data <= saw_rom(4054);
     when "111111010111" => data <= saw_rom(4055);
     when "111111011000" => data <= saw_rom(4056);
     when "111111011001" => data <= saw_rom(4057);
     when "111111011010" => data <= saw_rom(4058);
     when "111111011011" => data <= saw_rom(4059);
     when "111111011100" => data <= saw_rom(4060);
     when "111111011101" => data <= saw_rom(4061);
     when "111111011110" => data <= saw_rom(4062);
     when "111111011111" => data <= saw_rom(4063);
     when "111111100000" => data <= saw_rom(4064);
     when "111111100001" => data <= saw_rom(4065);
     when "111111100010" => data <= saw_rom(4066);
     when "111111100011" => data <= saw_rom(4067);
     when "111111100100" => data <= saw_rom(4068);
     when "111111100101" => data <= saw_rom(4069);
     when "111111100110" => data <= saw_rom(4070);
     when "111111100111" => data <= saw_rom(4071);
     when "111111101000" => data <= saw_rom(4072);
     when "111111101001" => data <= saw_rom(4073);
     when "111111101010" => data <= saw_rom(4074);
     when "111111101011" => data <= saw_rom(4075);
     when "111111101100" => data <= saw_rom(4076);
     when "111111101101" => data <= saw_rom(4077);
     when "111111101110" => data <= saw_rom(4078);
     when "111111101111" => data <= saw_rom(4079);
     when "111111110000" => data <= saw_rom(4080);
     when "111111110001" => data <= saw_rom(4081);
     when "111111110010" => data <= saw_rom(4082);
     when "111111110011" => data <= saw_rom(4083);
     when "111111110100" => data <= saw_rom(4084);
     when "111111110101" => data <= saw_rom(4085);
     when "111111110110" => data <= saw_rom(4086);
     when "111111110111" => data <= saw_rom(4087);
     when "111111111000" => data <= saw_rom(4088);
     when "111111111001" => data <= saw_rom(4089);
     when "111111111010" => data <= saw_rom(4090);
     when "111111111011" => data <= saw_rom(4091);
     when "111111111100" => data <= saw_rom(4092);
     when "111111111101" => data <= saw_rom(4093);
     when "111111111110" => data <= saw_rom(4094);
     when "111111111111" => data <= saw_rom(4095);
     when others => data <= "000000000000";
    end case;
 end process;
end arch_Sawtooth_LUT;
