library ieee;
use ieee.std_logic_1164.all;
entity Triangle_LUT is
 port ( address : in std_logic_vector(11 downto 0);
    data : out std_logic_vector(11 downto 0));
 end entity Triangle_LUT;
 architecture arch_Triangle_LUT of Triangle_LUT is
    type mem is array ( 0 to 2**12 - 1) of std_logic_vector(11 downto 0);
    constant triangle_rom : mem := (
    0 => "000000000000",
    1 => "000000000010",
    2 => "000000000100",
    3 => "000000000110",
    4 => "000000001000",
    5 => "000000001010",
    6 => "000000001100",
    7 => "000000001110",
    8 => "000000010000",
    9 => "000000010010",
    10 => "000000010100",
    11 => "000000010110",
    12 => "000000011000",
    13 => "000000011010",
    14 => "000000011100",
    15 => "000000011110",
    16 => "000000100000",
    17 => "000000100010",
    18 => "000000100100",
    19 => "000000100110",
    20 => "000000101000",
    21 => "000000101010",
    22 => "000000101100",
    23 => "000000101110",
    24 => "000000110000",
    25 => "000000110010",
    26 => "000000110100",
    27 => "000000110110",
    28 => "000000111000",
    29 => "000000111010",
    30 => "000000111100",
    31 => "000000111110",
    32 => "000001000000",
    33 => "000001000010",
    34 => "000001000100",
    35 => "000001000110",
    36 => "000001001000",
    37 => "000001001010",
    38 => "000001001100",
    39 => "000001001110",
    40 => "000001010000",
    41 => "000001010010",
    42 => "000001010100",
    43 => "000001010110",
    44 => "000001011000",
    45 => "000001011010",
    46 => "000001011100",
    47 => "000001011110",
    48 => "000001100000",
    49 => "000001100010",
    50 => "000001100100",
    51 => "000001100110",
    52 => "000001101000",
    53 => "000001101010",
    54 => "000001101100",
    55 => "000001101110",
    56 => "000001110000",
    57 => "000001110010",
    58 => "000001110100",
    59 => "000001110110",
    60 => "000001111000",
    61 => "000001111010",
    62 => "000001111100",
    63 => "000001111110",
    64 => "000010000000",
    65 => "000010000010",
    66 => "000010000100",
    67 => "000010000110",
    68 => "000010001000",
    69 => "000010001010",
    70 => "000010001100",
    71 => "000010001110",
    72 => "000010010000",
    73 => "000010010010",
    74 => "000010010100",
    75 => "000010010110",
    76 => "000010011000",
    77 => "000010011010",
    78 => "000010011100",
    79 => "000010011110",
    80 => "000010100000",
    81 => "000010100010",
    82 => "000010100100",
    83 => "000010100110",
    84 => "000010101000",
    85 => "000010101010",
    86 => "000010101100",
    87 => "000010101110",
    88 => "000010110000",
    89 => "000010110010",
    90 => "000010110100",
    91 => "000010110110",
    92 => "000010111000",
    93 => "000010111010",
    94 => "000010111100",
    95 => "000010111110",
    96 => "000011000000",
    97 => "000011000010",
    98 => "000011000100",
    99 => "000011000110",
    100 => "000011001000",
    101 => "000011001010",
    102 => "000011001100",
    103 => "000011001110",
    104 => "000011010000",
    105 => "000011010010",
    106 => "000011010100",
    107 => "000011010110",
    108 => "000011011000",
    109 => "000011011010",
    110 => "000011011100",
    111 => "000011011110",
    112 => "000011100000",
    113 => "000011100010",
    114 => "000011100100",
    115 => "000011100110",
    116 => "000011101000",
    117 => "000011101010",
    118 => "000011101100",
    119 => "000011101110",
    120 => "000011110000",
    121 => "000011110010",
    122 => "000011110100",
    123 => "000011110110",
    124 => "000011111000",
    125 => "000011111010",
    126 => "000011111100",
    127 => "000011111110",
    128 => "000100000000",
    129 => "000100000010",
    130 => "000100000100",
    131 => "000100000110",
    132 => "000100001000",
    133 => "000100001010",
    134 => "000100001100",
    135 => "000100001110",
    136 => "000100010000",
    137 => "000100010010",
    138 => "000100010100",
    139 => "000100010110",
    140 => "000100011000",
    141 => "000100011010",
    142 => "000100011100",
    143 => "000100011110",
    144 => "000100100000",
    145 => "000100100010",
    146 => "000100100100",
    147 => "000100100110",
    148 => "000100101000",
    149 => "000100101010",
    150 => "000100101100",
    151 => "000100101110",
    152 => "000100110000",
    153 => "000100110010",
    154 => "000100110100",
    155 => "000100110110",
    156 => "000100111000",
    157 => "000100111010",
    158 => "000100111100",
    159 => "000100111110",
    160 => "000101000000",
    161 => "000101000010",
    162 => "000101000100",
    163 => "000101000110",
    164 => "000101001000",
    165 => "000101001010",
    166 => "000101001100",
    167 => "000101001110",
    168 => "000101010000",
    169 => "000101010010",
    170 => "000101010100",
    171 => "000101010110",
    172 => "000101011000",
    173 => "000101011010",
    174 => "000101011100",
    175 => "000101011110",
    176 => "000101100000",
    177 => "000101100010",
    178 => "000101100100",
    179 => "000101100110",
    180 => "000101101000",
    181 => "000101101010",
    182 => "000101101100",
    183 => "000101101110",
    184 => "000101110000",
    185 => "000101110010",
    186 => "000101110100",
    187 => "000101110110",
    188 => "000101111000",
    189 => "000101111010",
    190 => "000101111100",
    191 => "000101111110",
    192 => "000110000000",
    193 => "000110000010",
    194 => "000110000100",
    195 => "000110000110",
    196 => "000110001000",
    197 => "000110001010",
    198 => "000110001100",
    199 => "000110001110",
    200 => "000110010000",
    201 => "000110010010",
    202 => "000110010100",
    203 => "000110010110",
    204 => "000110011000",
    205 => "000110011010",
    206 => "000110011100",
    207 => "000110011110",
    208 => "000110100000",
    209 => "000110100010",
    210 => "000110100100",
    211 => "000110100110",
    212 => "000110101000",
    213 => "000110101010",
    214 => "000110101100",
    215 => "000110101110",
    216 => "000110110000",
    217 => "000110110010",
    218 => "000110110100",
    219 => "000110110110",
    220 => "000110111000",
    221 => "000110111010",
    222 => "000110111100",
    223 => "000110111110",
    224 => "000111000000",
    225 => "000111000010",
    226 => "000111000100",
    227 => "000111000110",
    228 => "000111001000",
    229 => "000111001010",
    230 => "000111001100",
    231 => "000111001110",
    232 => "000111010000",
    233 => "000111010010",
    234 => "000111010100",
    235 => "000111010110",
    236 => "000111011000",
    237 => "000111011010",
    238 => "000111011100",
    239 => "000111011110",
    240 => "000111100000",
    241 => "000111100010",
    242 => "000111100100",
    243 => "000111100110",
    244 => "000111101000",
    245 => "000111101010",
    246 => "000111101100",
    247 => "000111101110",
    248 => "000111110000",
    249 => "000111110010",
    250 => "000111110100",
    251 => "000111110110",
    252 => "000111111000",
    253 => "000111111010",
    254 => "000111111100",
    255 => "000111111110",
    256 => "001000000000",
    257 => "001000000010",
    258 => "001000000100",
    259 => "001000000110",
    260 => "001000001000",
    261 => "001000001010",
    262 => "001000001100",
    263 => "001000001110",
    264 => "001000010000",
    265 => "001000010010",
    266 => "001000010100",
    267 => "001000010110",
    268 => "001000011000",
    269 => "001000011010",
    270 => "001000011100",
    271 => "001000011110",
    272 => "001000100000",
    273 => "001000100010",
    274 => "001000100100",
    275 => "001000100110",
    276 => "001000101000",
    277 => "001000101010",
    278 => "001000101100",
    279 => "001000101110",
    280 => "001000110000",
    281 => "001000110010",
    282 => "001000110100",
    283 => "001000110110",
    284 => "001000111000",
    285 => "001000111010",
    286 => "001000111100",
    287 => "001000111110",
    288 => "001001000000",
    289 => "001001000010",
    290 => "001001000100",
    291 => "001001000110",
    292 => "001001001000",
    293 => "001001001010",
    294 => "001001001100",
    295 => "001001001110",
    296 => "001001010000",
    297 => "001001010010",
    298 => "001001010100",
    299 => "001001010110",
    300 => "001001011000",
    301 => "001001011010",
    302 => "001001011100",
    303 => "001001011110",
    304 => "001001100000",
    305 => "001001100010",
    306 => "001001100100",
    307 => "001001100110",
    308 => "001001101000",
    309 => "001001101010",
    310 => "001001101100",
    311 => "001001101110",
    312 => "001001110000",
    313 => "001001110010",
    314 => "001001110100",
    315 => "001001110110",
    316 => "001001111000",
    317 => "001001111010",
    318 => "001001111100",
    319 => "001001111110",
    320 => "001010000000",
    321 => "001010000010",
    322 => "001010000100",
    323 => "001010000110",
    324 => "001010001000",
    325 => "001010001010",
    326 => "001010001100",
    327 => "001010001110",
    328 => "001010010000",
    329 => "001010010010",
    330 => "001010010100",
    331 => "001010010110",
    332 => "001010011000",
    333 => "001010011010",
    334 => "001010011100",
    335 => "001010011110",
    336 => "001010100000",
    337 => "001010100010",
    338 => "001010100100",
    339 => "001010100110",
    340 => "001010101000",
    341 => "001010101010",
    342 => "001010101100",
    343 => "001010101110",
    344 => "001010110000",
    345 => "001010110010",
    346 => "001010110100",
    347 => "001010110110",
    348 => "001010111000",
    349 => "001010111010",
    350 => "001010111100",
    351 => "001010111110",
    352 => "001011000000",
    353 => "001011000010",
    354 => "001011000100",
    355 => "001011000110",
    356 => "001011001000",
    357 => "001011001010",
    358 => "001011001100",
    359 => "001011001110",
    360 => "001011010000",
    361 => "001011010010",
    362 => "001011010100",
    363 => "001011010110",
    364 => "001011011000",
    365 => "001011011010",
    366 => "001011011100",
    367 => "001011011110",
    368 => "001011100000",
    369 => "001011100010",
    370 => "001011100100",
    371 => "001011100110",
    372 => "001011101000",
    373 => "001011101010",
    374 => "001011101100",
    375 => "001011101110",
    376 => "001011110000",
    377 => "001011110010",
    378 => "001011110100",
    379 => "001011110110",
    380 => "001011111000",
    381 => "001011111010",
    382 => "001011111100",
    383 => "001011111110",
    384 => "001100000000",
    385 => "001100000010",
    386 => "001100000100",
    387 => "001100000110",
    388 => "001100001000",
    389 => "001100001010",
    390 => "001100001100",
    391 => "001100001110",
    392 => "001100010000",
    393 => "001100010010",
    394 => "001100010100",
    395 => "001100010110",
    396 => "001100011000",
    397 => "001100011010",
    398 => "001100011100",
    399 => "001100011110",
    400 => "001100100000",
    401 => "001100100010",
    402 => "001100100100",
    403 => "001100100110",
    404 => "001100101000",
    405 => "001100101010",
    406 => "001100101100",
    407 => "001100101110",
    408 => "001100110000",
    409 => "001100110010",
    410 => "001100110100",
    411 => "001100110110",
    412 => "001100111000",
    413 => "001100111010",
    414 => "001100111100",
    415 => "001100111110",
    416 => "001101000000",
    417 => "001101000010",
    418 => "001101000100",
    419 => "001101000110",
    420 => "001101001000",
    421 => "001101001010",
    422 => "001101001100",
    423 => "001101001110",
    424 => "001101010000",
    425 => "001101010010",
    426 => "001101010100",
    427 => "001101010110",
    428 => "001101011000",
    429 => "001101011010",
    430 => "001101011100",
    431 => "001101011110",
    432 => "001101100000",
    433 => "001101100010",
    434 => "001101100100",
    435 => "001101100110",
    436 => "001101101000",
    437 => "001101101010",
    438 => "001101101100",
    439 => "001101101110",
    440 => "001101110000",
    441 => "001101110010",
    442 => "001101110100",
    443 => "001101110110",
    444 => "001101111000",
    445 => "001101111010",
    446 => "001101111100",
    447 => "001101111110",
    448 => "001110000000",
    449 => "001110000010",
    450 => "001110000100",
    451 => "001110000110",
    452 => "001110001000",
    453 => "001110001010",
    454 => "001110001100",
    455 => "001110001110",
    456 => "001110010000",
    457 => "001110010010",
    458 => "001110010100",
    459 => "001110010110",
    460 => "001110011000",
    461 => "001110011010",
    462 => "001110011100",
    463 => "001110011110",
    464 => "001110100000",
    465 => "001110100010",
    466 => "001110100100",
    467 => "001110100110",
    468 => "001110101000",
    469 => "001110101010",
    470 => "001110101100",
    471 => "001110101110",
    472 => "001110110000",
    473 => "001110110010",
    474 => "001110110100",
    475 => "001110110110",
    476 => "001110111000",
    477 => "001110111010",
    478 => "001110111100",
    479 => "001110111110",
    480 => "001111000000",
    481 => "001111000010",
    482 => "001111000100",
    483 => "001111000110",
    484 => "001111001000",
    485 => "001111001010",
    486 => "001111001100",
    487 => "001111001110",
    488 => "001111010000",
    489 => "001111010010",
    490 => "001111010100",
    491 => "001111010110",
    492 => "001111011000",
    493 => "001111011010",
    494 => "001111011100",
    495 => "001111011110",
    496 => "001111100000",
    497 => "001111100010",
    498 => "001111100100",
    499 => "001111100110",
    500 => "001111101000",
    501 => "001111101010",
    502 => "001111101100",
    503 => "001111101110",
    504 => "001111110000",
    505 => "001111110010",
    506 => "001111110100",
    507 => "001111110110",
    508 => "001111111000",
    509 => "001111111010",
    510 => "001111111100",
    511 => "001111111110",
    512 => "010000000000",
    513 => "010000000010",
    514 => "010000000100",
    515 => "010000000110",
    516 => "010000001000",
    517 => "010000001010",
    518 => "010000001100",
    519 => "010000001110",
    520 => "010000010000",
    521 => "010000010010",
    522 => "010000010100",
    523 => "010000010110",
    524 => "010000011000",
    525 => "010000011010",
    526 => "010000011100",
    527 => "010000011110",
    528 => "010000100000",
    529 => "010000100010",
    530 => "010000100100",
    531 => "010000100110",
    532 => "010000101000",
    533 => "010000101010",
    534 => "010000101100",
    535 => "010000101110",
    536 => "010000110000",
    537 => "010000110010",
    538 => "010000110100",
    539 => "010000110110",
    540 => "010000111000",
    541 => "010000111010",
    542 => "010000111100",
    543 => "010000111110",
    544 => "010001000000",
    545 => "010001000010",
    546 => "010001000100",
    547 => "010001000110",
    548 => "010001001000",
    549 => "010001001010",
    550 => "010001001100",
    551 => "010001001110",
    552 => "010001010000",
    553 => "010001010010",
    554 => "010001010100",
    555 => "010001010110",
    556 => "010001011000",
    557 => "010001011010",
    558 => "010001011100",
    559 => "010001011110",
    560 => "010001100000",
    561 => "010001100010",
    562 => "010001100100",
    563 => "010001100110",
    564 => "010001101000",
    565 => "010001101010",
    566 => "010001101100",
    567 => "010001101110",
    568 => "010001110000",
    569 => "010001110010",
    570 => "010001110100",
    571 => "010001110110",
    572 => "010001111000",
    573 => "010001111010",
    574 => "010001111100",
    575 => "010001111110",
    576 => "010010000000",
    577 => "010010000010",
    578 => "010010000100",
    579 => "010010000110",
    580 => "010010001000",
    581 => "010010001010",
    582 => "010010001100",
    583 => "010010001110",
    584 => "010010010000",
    585 => "010010010010",
    586 => "010010010100",
    587 => "010010010110",
    588 => "010010011000",
    589 => "010010011010",
    590 => "010010011100",
    591 => "010010011110",
    592 => "010010100000",
    593 => "010010100010",
    594 => "010010100100",
    595 => "010010100110",
    596 => "010010101000",
    597 => "010010101010",
    598 => "010010101100",
    599 => "010010101110",
    600 => "010010110000",
    601 => "010010110010",
    602 => "010010110100",
    603 => "010010110110",
    604 => "010010111000",
    605 => "010010111010",
    606 => "010010111100",
    607 => "010010111110",
    608 => "010011000000",
    609 => "010011000010",
    610 => "010011000100",
    611 => "010011000110",
    612 => "010011001000",
    613 => "010011001010",
    614 => "010011001100",
    615 => "010011001110",
    616 => "010011010000",
    617 => "010011010010",
    618 => "010011010100",
    619 => "010011010110",
    620 => "010011011000",
    621 => "010011011010",
    622 => "010011011100",
    623 => "010011011110",
    624 => "010011100000",
    625 => "010011100010",
    626 => "010011100100",
    627 => "010011100110",
    628 => "010011101000",
    629 => "010011101010",
    630 => "010011101100",
    631 => "010011101110",
    632 => "010011110000",
    633 => "010011110010",
    634 => "010011110100",
    635 => "010011110110",
    636 => "010011111000",
    637 => "010011111010",
    638 => "010011111100",
    639 => "010011111110",
    640 => "010100000000",
    641 => "010100000010",
    642 => "010100000100",
    643 => "010100000110",
    644 => "010100001000",
    645 => "010100001010",
    646 => "010100001100",
    647 => "010100001110",
    648 => "010100010000",
    649 => "010100010010",
    650 => "010100010100",
    651 => "010100010110",
    652 => "010100011000",
    653 => "010100011010",
    654 => "010100011100",
    655 => "010100011110",
    656 => "010100100000",
    657 => "010100100010",
    658 => "010100100100",
    659 => "010100100110",
    660 => "010100101000",
    661 => "010100101010",
    662 => "010100101100",
    663 => "010100101110",
    664 => "010100110000",
    665 => "010100110010",
    666 => "010100110100",
    667 => "010100110110",
    668 => "010100111000",
    669 => "010100111010",
    670 => "010100111100",
    671 => "010100111110",
    672 => "010101000000",
    673 => "010101000010",
    674 => "010101000100",
    675 => "010101000110",
    676 => "010101001000",
    677 => "010101001010",
    678 => "010101001100",
    679 => "010101001110",
    680 => "010101010000",
    681 => "010101010010",
    682 => "010101010100",
    683 => "010101010110",
    684 => "010101011000",
    685 => "010101011010",
    686 => "010101011100",
    687 => "010101011110",
    688 => "010101100000",
    689 => "010101100010",
    690 => "010101100100",
    691 => "010101100110",
    692 => "010101101000",
    693 => "010101101010",
    694 => "010101101100",
    695 => "010101101110",
    696 => "010101110000",
    697 => "010101110010",
    698 => "010101110100",
    699 => "010101110110",
    700 => "010101111000",
    701 => "010101111010",
    702 => "010101111100",
    703 => "010101111110",
    704 => "010110000000",
    705 => "010110000010",
    706 => "010110000100",
    707 => "010110000110",
    708 => "010110001000",
    709 => "010110001010",
    710 => "010110001100",
    711 => "010110001110",
    712 => "010110010000",
    713 => "010110010010",
    714 => "010110010100",
    715 => "010110010110",
    716 => "010110011000",
    717 => "010110011010",
    718 => "010110011100",
    719 => "010110011110",
    720 => "010110100000",
    721 => "010110100010",
    722 => "010110100100",
    723 => "010110100110",
    724 => "010110101000",
    725 => "010110101010",
    726 => "010110101100",
    727 => "010110101110",
    728 => "010110110000",
    729 => "010110110010",
    730 => "010110110100",
    731 => "010110110110",
    732 => "010110111000",
    733 => "010110111010",
    734 => "010110111100",
    735 => "010110111110",
    736 => "010111000000",
    737 => "010111000010",
    738 => "010111000100",
    739 => "010111000110",
    740 => "010111001000",
    741 => "010111001010",
    742 => "010111001100",
    743 => "010111001110",
    744 => "010111010000",
    745 => "010111010010",
    746 => "010111010100",
    747 => "010111010110",
    748 => "010111011000",
    749 => "010111011010",
    750 => "010111011100",
    751 => "010111011110",
    752 => "010111100000",
    753 => "010111100010",
    754 => "010111100100",
    755 => "010111100110",
    756 => "010111101000",
    757 => "010111101010",
    758 => "010111101100",
    759 => "010111101110",
    760 => "010111110000",
    761 => "010111110010",
    762 => "010111110100",
    763 => "010111110110",
    764 => "010111111000",
    765 => "010111111010",
    766 => "010111111100",
    767 => "010111111110",
    768 => "011000000000",
    769 => "011000000010",
    770 => "011000000100",
    771 => "011000000110",
    772 => "011000001000",
    773 => "011000001010",
    774 => "011000001100",
    775 => "011000001110",
    776 => "011000010000",
    777 => "011000010010",
    778 => "011000010100",
    779 => "011000010110",
    780 => "011000011000",
    781 => "011000011010",
    782 => "011000011100",
    783 => "011000011110",
    784 => "011000100000",
    785 => "011000100010",
    786 => "011000100100",
    787 => "011000100110",
    788 => "011000101000",
    789 => "011000101010",
    790 => "011000101100",
    791 => "011000101110",
    792 => "011000110000",
    793 => "011000110010",
    794 => "011000110100",
    795 => "011000110110",
    796 => "011000111000",
    797 => "011000111010",
    798 => "011000111100",
    799 => "011000111110",
    800 => "011001000000",
    801 => "011001000010",
    802 => "011001000100",
    803 => "011001000110",
    804 => "011001001000",
    805 => "011001001010",
    806 => "011001001100",
    807 => "011001001110",
    808 => "011001010000",
    809 => "011001010010",
    810 => "011001010100",
    811 => "011001010110",
    812 => "011001011000",
    813 => "011001011010",
    814 => "011001011100",
    815 => "011001011110",
    816 => "011001100000",
    817 => "011001100010",
    818 => "011001100100",
    819 => "011001100110",
    820 => "011001101000",
    821 => "011001101010",
    822 => "011001101100",
    823 => "011001101110",
    824 => "011001110000",
    825 => "011001110010",
    826 => "011001110100",
    827 => "011001110110",
    828 => "011001111000",
    829 => "011001111010",
    830 => "011001111100",
    831 => "011001111110",
    832 => "011010000000",
    833 => "011010000010",
    834 => "011010000011",
    835 => "011010000101",
    836 => "011010000111",
    837 => "011010001001",
    838 => "011010001011",
    839 => "011010001101",
    840 => "011010001111",
    841 => "011010010001",
    842 => "011010010011",
    843 => "011010010101",
    844 => "011010010111",
    845 => "011010011001",
    846 => "011010011011",
    847 => "011010011101",
    848 => "011010011111",
    849 => "011010100001",
    850 => "011010100011",
    851 => "011010100101",
    852 => "011010100111",
    853 => "011010101001",
    854 => "011010101011",
    855 => "011010101101",
    856 => "011010101111",
    857 => "011010110001",
    858 => "011010110011",
    859 => "011010110101",
    860 => "011010110111",
    861 => "011010111001",
    862 => "011010111011",
    863 => "011010111101",
    864 => "011010111111",
    865 => "011011000001",
    866 => "011011000011",
    867 => "011011000101",
    868 => "011011000111",
    869 => "011011001001",
    870 => "011011001011",
    871 => "011011001101",
    872 => "011011001111",
    873 => "011011010001",
    874 => "011011010011",
    875 => "011011010101",
    876 => "011011010111",
    877 => "011011011001",
    878 => "011011011011",
    879 => "011011011101",
    880 => "011011011111",
    881 => "011011100001",
    882 => "011011100011",
    883 => "011011100101",
    884 => "011011100111",
    885 => "011011101001",
    886 => "011011101011",
    887 => "011011101101",
    888 => "011011101111",
    889 => "011011110001",
    890 => "011011110011",
    891 => "011011110101",
    892 => "011011110111",
    893 => "011011111001",
    894 => "011011111011",
    895 => "011011111101",
    896 => "011011111111",
    897 => "011100000001",
    898 => "011100000011",
    899 => "011100000101",
    900 => "011100000111",
    901 => "011100001001",
    902 => "011100001011",
    903 => "011100001101",
    904 => "011100001111",
    905 => "011100010001",
    906 => "011100010011",
    907 => "011100010101",
    908 => "011100010111",
    909 => "011100011001",
    910 => "011100011011",
    911 => "011100011101",
    912 => "011100011111",
    913 => "011100100001",
    914 => "011100100011",
    915 => "011100100101",
    916 => "011100100111",
    917 => "011100101001",
    918 => "011100101011",
    919 => "011100101101",
    920 => "011100101111",
    921 => "011100110001",
    922 => "011100110011",
    923 => "011100110101",
    924 => "011100110111",
    925 => "011100111001",
    926 => "011100111011",
    927 => "011100111101",
    928 => "011100111111",
    929 => "011101000001",
    930 => "011101000011",
    931 => "011101000101",
    932 => "011101000111",
    933 => "011101001001",
    934 => "011101001011",
    935 => "011101001101",
    936 => "011101001111",
    937 => "011101010001",
    938 => "011101010011",
    939 => "011101010101",
    940 => "011101010111",
    941 => "011101011001",
    942 => "011101011011",
    943 => "011101011101",
    944 => "011101011111",
    945 => "011101100001",
    946 => "011101100011",
    947 => "011101100101",
    948 => "011101100111",
    949 => "011101101001",
    950 => "011101101011",
    951 => "011101101101",
    952 => "011101101111",
    953 => "011101110001",
    954 => "011101110011",
    955 => "011101110101",
    956 => "011101110111",
    957 => "011101111001",
    958 => "011101111011",
    959 => "011101111101",
    960 => "011101111111",
    961 => "011110000001",
    962 => "011110000011",
    963 => "011110000101",
    964 => "011110000111",
    965 => "011110001001",
    966 => "011110001011",
    967 => "011110001101",
    968 => "011110001111",
    969 => "011110010001",
    970 => "011110010011",
    971 => "011110010101",
    972 => "011110010111",
    973 => "011110011001",
    974 => "011110011011",
    975 => "011110011101",
    976 => "011110011111",
    977 => "011110100001",
    978 => "011110100011",
    979 => "011110100101",
    980 => "011110100111",
    981 => "011110101001",
    982 => "011110101011",
    983 => "011110101101",
    984 => "011110101111",
    985 => "011110110001",
    986 => "011110110011",
    987 => "011110110101",
    988 => "011110110111",
    989 => "011110111001",
    990 => "011110111011",
    991 => "011110111101",
    992 => "011110111111",
    993 => "011111000001",
    994 => "011111000011",
    995 => "011111000101",
    996 => "011111000111",
    997 => "011111001001",
    998 => "011111001011",
    999 => "011111001101",
    1000 => "011111001111",
    1001 => "011111010001",
    1002 => "011111010011",
    1003 => "011111010101",
    1004 => "011111010111",
    1005 => "011111011001",
    1006 => "011111011011",
    1007 => "011111011101",
    1008 => "011111011111",
    1009 => "011111100001",
    1010 => "011111100011",
    1011 => "011111100101",
    1012 => "011111100111",
    1013 => "011111101001",
    1014 => "011111101011",
    1015 => "011111101101",
    1016 => "011111101111",
    1017 => "011111110001",
    1018 => "011111110011",
    1019 => "011111110101",
    1020 => "011111110111",
    1021 => "011111111001",
    1022 => "011111111011",
    1023 => "011111111101",
    1024 => "011111111111",
    1025 => "100000000001",
    1026 => "100000000011",
    1027 => "100000000101",
    1028 => "100000000111",
    1029 => "100000001001",
    1030 => "100000001011",
    1031 => "100000001101",
    1032 => "100000001111",
    1033 => "100000010001",
    1034 => "100000010011",
    1035 => "100000010101",
    1036 => "100000010111",
    1037 => "100000011001",
    1038 => "100000011011",
    1039 => "100000011101",
    1040 => "100000011111",
    1041 => "100000100001",
    1042 => "100000100011",
    1043 => "100000100101",
    1044 => "100000100111",
    1045 => "100000101001",
    1046 => "100000101011",
    1047 => "100000101101",
    1048 => "100000101111",
    1049 => "100000110001",
    1050 => "100000110011",
    1051 => "100000110101",
    1052 => "100000110111",
    1053 => "100000111001",
    1054 => "100000111011",
    1055 => "100000111101",
    1056 => "100000111111",
    1057 => "100001000001",
    1058 => "100001000011",
    1059 => "100001000101",
    1060 => "100001000111",
    1061 => "100001001001",
    1062 => "100001001011",
    1063 => "100001001101",
    1064 => "100001001111",
    1065 => "100001010001",
    1066 => "100001010011",
    1067 => "100001010101",
    1068 => "100001010111",
    1069 => "100001011001",
    1070 => "100001011011",
    1071 => "100001011101",
    1072 => "100001011111",
    1073 => "100001100001",
    1074 => "100001100011",
    1075 => "100001100101",
    1076 => "100001100111",
    1077 => "100001101001",
    1078 => "100001101011",
    1079 => "100001101101",
    1080 => "100001101111",
    1081 => "100001110001",
    1082 => "100001110011",
    1083 => "100001110101",
    1084 => "100001110111",
    1085 => "100001111001",
    1086 => "100001111011",
    1087 => "100001111101",
    1088 => "100001111111",
    1089 => "100010000001",
    1090 => "100010000011",
    1091 => "100010000101",
    1092 => "100010000111",
    1093 => "100010001001",
    1094 => "100010001011",
    1095 => "100010001101",
    1096 => "100010001111",
    1097 => "100010010001",
    1098 => "100010010011",
    1099 => "100010010101",
    1100 => "100010010111",
    1101 => "100010011001",
    1102 => "100010011011",
    1103 => "100010011101",
    1104 => "100010011111",
    1105 => "100010100001",
    1106 => "100010100011",
    1107 => "100010100101",
    1108 => "100010100111",
    1109 => "100010101001",
    1110 => "100010101011",
    1111 => "100010101101",
    1112 => "100010101111",
    1113 => "100010110001",
    1114 => "100010110011",
    1115 => "100010110101",
    1116 => "100010110111",
    1117 => "100010111001",
    1118 => "100010111011",
    1119 => "100010111101",
    1120 => "100010111111",
    1121 => "100011000001",
    1122 => "100011000011",
    1123 => "100011000101",
    1124 => "100011000111",
    1125 => "100011001001",
    1126 => "100011001011",
    1127 => "100011001101",
    1128 => "100011001111",
    1129 => "100011010001",
    1130 => "100011010011",
    1131 => "100011010101",
    1132 => "100011010111",
    1133 => "100011011001",
    1134 => "100011011011",
    1135 => "100011011101",
    1136 => "100011011111",
    1137 => "100011100001",
    1138 => "100011100011",
    1139 => "100011100101",
    1140 => "100011100111",
    1141 => "100011101001",
    1142 => "100011101011",
    1143 => "100011101101",
    1144 => "100011101111",
    1145 => "100011110001",
    1146 => "100011110011",
    1147 => "100011110101",
    1148 => "100011110111",
    1149 => "100011111001",
    1150 => "100011111011",
    1151 => "100011111101",
    1152 => "100011111111",
    1153 => "100100000001",
    1154 => "100100000011",
    1155 => "100100000101",
    1156 => "100100000111",
    1157 => "100100001001",
    1158 => "100100001011",
    1159 => "100100001101",
    1160 => "100100001111",
    1161 => "100100010001",
    1162 => "100100010011",
    1163 => "100100010101",
    1164 => "100100010111",
    1165 => "100100011001",
    1166 => "100100011011",
    1167 => "100100011101",
    1168 => "100100011111",
    1169 => "100100100001",
    1170 => "100100100011",
    1171 => "100100100101",
    1172 => "100100100111",
    1173 => "100100101001",
    1174 => "100100101011",
    1175 => "100100101101",
    1176 => "100100101111",
    1177 => "100100110001",
    1178 => "100100110011",
    1179 => "100100110101",
    1180 => "100100110111",
    1181 => "100100111001",
    1182 => "100100111011",
    1183 => "100100111101",
    1184 => "100100111111",
    1185 => "100101000001",
    1186 => "100101000011",
    1187 => "100101000101",
    1188 => "100101000111",
    1189 => "100101001001",
    1190 => "100101001011",
    1191 => "100101001101",
    1192 => "100101001111",
    1193 => "100101010001",
    1194 => "100101010011",
    1195 => "100101010101",
    1196 => "100101010111",
    1197 => "100101011001",
    1198 => "100101011011",
    1199 => "100101011101",
    1200 => "100101011111",
    1201 => "100101100001",
    1202 => "100101100011",
    1203 => "100101100101",
    1204 => "100101100111",
    1205 => "100101101001",
    1206 => "100101101011",
    1207 => "100101101101",
    1208 => "100101101111",
    1209 => "100101110001",
    1210 => "100101110011",
    1211 => "100101110101",
    1212 => "100101110111",
    1213 => "100101111001",
    1214 => "100101111011",
    1215 => "100101111101",
    1216 => "100101111111",
    1217 => "100110000001",
    1218 => "100110000011",
    1219 => "100110000101",
    1220 => "100110000111",
    1221 => "100110001001",
    1222 => "100110001011",
    1223 => "100110001101",
    1224 => "100110001111",
    1225 => "100110010001",
    1226 => "100110010011",
    1227 => "100110010101",
    1228 => "100110010111",
    1229 => "100110011001",
    1230 => "100110011011",
    1231 => "100110011101",
    1232 => "100110011111",
    1233 => "100110100001",
    1234 => "100110100011",
    1235 => "100110100101",
    1236 => "100110100111",
    1237 => "100110101001",
    1238 => "100110101011",
    1239 => "100110101101",
    1240 => "100110101111",
    1241 => "100110110001",
    1242 => "100110110011",
    1243 => "100110110101",
    1244 => "100110110111",
    1245 => "100110111001",
    1246 => "100110111011",
    1247 => "100110111101",
    1248 => "100110111111",
    1249 => "100111000001",
    1250 => "100111000011",
    1251 => "100111000101",
    1252 => "100111000111",
    1253 => "100111001001",
    1254 => "100111001011",
    1255 => "100111001101",
    1256 => "100111001111",
    1257 => "100111010001",
    1258 => "100111010011",
    1259 => "100111010101",
    1260 => "100111010111",
    1261 => "100111011001",
    1262 => "100111011011",
    1263 => "100111011101",
    1264 => "100111011111",
    1265 => "100111100001",
    1266 => "100111100011",
    1267 => "100111100101",
    1268 => "100111100111",
    1269 => "100111101001",
    1270 => "100111101011",
    1271 => "100111101101",
    1272 => "100111101111",
    1273 => "100111110001",
    1274 => "100111110011",
    1275 => "100111110101",
    1276 => "100111110111",
    1277 => "100111111001",
    1278 => "100111111011",
    1279 => "100111111101",
    1280 => "100111111111",
    1281 => "101000000001",
    1282 => "101000000011",
    1283 => "101000000101",
    1284 => "101000000111",
    1285 => "101000001001",
    1286 => "101000001011",
    1287 => "101000001101",
    1288 => "101000001111",
    1289 => "101000010001",
    1290 => "101000010011",
    1291 => "101000010101",
    1292 => "101000010111",
    1293 => "101000011001",
    1294 => "101000011011",
    1295 => "101000011101",
    1296 => "101000011111",
    1297 => "101000100001",
    1298 => "101000100011",
    1299 => "101000100101",
    1300 => "101000100111",
    1301 => "101000101001",
    1302 => "101000101011",
    1303 => "101000101101",
    1304 => "101000101111",
    1305 => "101000110001",
    1306 => "101000110011",
    1307 => "101000110101",
    1308 => "101000110111",
    1309 => "101000111001",
    1310 => "101000111011",
    1311 => "101000111101",
    1312 => "101000111111",
    1313 => "101001000001",
    1314 => "101001000011",
    1315 => "101001000101",
    1316 => "101001000111",
    1317 => "101001001001",
    1318 => "101001001011",
    1319 => "101001001101",
    1320 => "101001001111",
    1321 => "101001010001",
    1322 => "101001010011",
    1323 => "101001010101",
    1324 => "101001010111",
    1325 => "101001011001",
    1326 => "101001011011",
    1327 => "101001011101",
    1328 => "101001011111",
    1329 => "101001100001",
    1330 => "101001100011",
    1331 => "101001100101",
    1332 => "101001100111",
    1333 => "101001101001",
    1334 => "101001101011",
    1335 => "101001101101",
    1336 => "101001101111",
    1337 => "101001110001",
    1338 => "101001110011",
    1339 => "101001110101",
    1340 => "101001110111",
    1341 => "101001111001",
    1342 => "101001111011",
    1343 => "101001111101",
    1344 => "101001111111",
    1345 => "101010000001",
    1346 => "101010000011",
    1347 => "101010000101",
    1348 => "101010000111",
    1349 => "101010001001",
    1350 => "101010001011",
    1351 => "101010001101",
    1352 => "101010001111",
    1353 => "101010010001",
    1354 => "101010010011",
    1355 => "101010010101",
    1356 => "101010010111",
    1357 => "101010011001",
    1358 => "101010011011",
    1359 => "101010011101",
    1360 => "101010011111",
    1361 => "101010100001",
    1362 => "101010100011",
    1363 => "101010100101",
    1364 => "101010100111",
    1365 => "101010101001",
    1366 => "101010101011",
    1367 => "101010101101",
    1368 => "101010101111",
    1369 => "101010110001",
    1370 => "101010110011",
    1371 => "101010110101",
    1372 => "101010110111",
    1373 => "101010111001",
    1374 => "101010111011",
    1375 => "101010111101",
    1376 => "101010111111",
    1377 => "101011000001",
    1378 => "101011000011",
    1379 => "101011000101",
    1380 => "101011000111",
    1381 => "101011001001",
    1382 => "101011001011",
    1383 => "101011001101",
    1384 => "101011001111",
    1385 => "101011010001",
    1386 => "101011010011",
    1387 => "101011010101",
    1388 => "101011010111",
    1389 => "101011011001",
    1390 => "101011011011",
    1391 => "101011011101",
    1392 => "101011011111",
    1393 => "101011100001",
    1394 => "101011100011",
    1395 => "101011100101",
    1396 => "101011100111",
    1397 => "101011101001",
    1398 => "101011101011",
    1399 => "101011101101",
    1400 => "101011101111",
    1401 => "101011110001",
    1402 => "101011110011",
    1403 => "101011110101",
    1404 => "101011110111",
    1405 => "101011111001",
    1406 => "101011111011",
    1407 => "101011111101",
    1408 => "101011111111",
    1409 => "101100000001",
    1410 => "101100000011",
    1411 => "101100000101",
    1412 => "101100000111",
    1413 => "101100001001",
    1414 => "101100001011",
    1415 => "101100001101",
    1416 => "101100001111",
    1417 => "101100010001",
    1418 => "101100010011",
    1419 => "101100010101",
    1420 => "101100010111",
    1421 => "101100011001",
    1422 => "101100011011",
    1423 => "101100011101",
    1424 => "101100011111",
    1425 => "101100100001",
    1426 => "101100100011",
    1427 => "101100100101",
    1428 => "101100100111",
    1429 => "101100101001",
    1430 => "101100101011",
    1431 => "101100101101",
    1432 => "101100101111",
    1433 => "101100110001",
    1434 => "101100110011",
    1435 => "101100110101",
    1436 => "101100110111",
    1437 => "101100111001",
    1438 => "101100111011",
    1439 => "101100111101",
    1440 => "101100111111",
    1441 => "101101000001",
    1442 => "101101000011",
    1443 => "101101000101",
    1444 => "101101000111",
    1445 => "101101001001",
    1446 => "101101001011",
    1447 => "101101001101",
    1448 => "101101001111",
    1449 => "101101010001",
    1450 => "101101010011",
    1451 => "101101010101",
    1452 => "101101010111",
    1453 => "101101011001",
    1454 => "101101011011",
    1455 => "101101011101",
    1456 => "101101011111",
    1457 => "101101100001",
    1458 => "101101100011",
    1459 => "101101100101",
    1460 => "101101100111",
    1461 => "101101101001",
    1462 => "101101101011",
    1463 => "101101101101",
    1464 => "101101101111",
    1465 => "101101110001",
    1466 => "101101110011",
    1467 => "101101110101",
    1468 => "101101110111",
    1469 => "101101111001",
    1470 => "101101111011",
    1471 => "101101111101",
    1472 => "101101111111",
    1473 => "101110000001",
    1474 => "101110000011",
    1475 => "101110000101",
    1476 => "101110000111",
    1477 => "101110001001",
    1478 => "101110001011",
    1479 => "101110001101",
    1480 => "101110001111",
    1481 => "101110010001",
    1482 => "101110010011",
    1483 => "101110010101",
    1484 => "101110010111",
    1485 => "101110011001",
    1486 => "101110011011",
    1487 => "101110011101",
    1488 => "101110011111",
    1489 => "101110100001",
    1490 => "101110100011",
    1491 => "101110100101",
    1492 => "101110100111",
    1493 => "101110101001",
    1494 => "101110101011",
    1495 => "101110101101",
    1496 => "101110101111",
    1497 => "101110110001",
    1498 => "101110110011",
    1499 => "101110110101",
    1500 => "101110110111",
    1501 => "101110111001",
    1502 => "101110111011",
    1503 => "101110111101",
    1504 => "101110111111",
    1505 => "101111000001",
    1506 => "101111000011",
    1507 => "101111000101",
    1508 => "101111000111",
    1509 => "101111001001",
    1510 => "101111001011",
    1511 => "101111001101",
    1512 => "101111001111",
    1513 => "101111010001",
    1514 => "101111010011",
    1515 => "101111010101",
    1516 => "101111010111",
    1517 => "101111011001",
    1518 => "101111011011",
    1519 => "101111011101",
    1520 => "101111011111",
    1521 => "101111100001",
    1522 => "101111100011",
    1523 => "101111100101",
    1524 => "101111100111",
    1525 => "101111101001",
    1526 => "101111101011",
    1527 => "101111101101",
    1528 => "101111101111",
    1529 => "101111110001",
    1530 => "101111110011",
    1531 => "101111110101",
    1532 => "101111110111",
    1533 => "101111111001",
    1534 => "101111111011",
    1535 => "101111111101",
    1536 => "101111111111",
    1537 => "110000000001",
    1538 => "110000000011",
    1539 => "110000000101",
    1540 => "110000000111",
    1541 => "110000001001",
    1542 => "110000001011",
    1543 => "110000001101",
    1544 => "110000001111",
    1545 => "110000010001",
    1546 => "110000010011",
    1547 => "110000010101",
    1548 => "110000010111",
    1549 => "110000011001",
    1550 => "110000011011",
    1551 => "110000011101",
    1552 => "110000011111",
    1553 => "110000100001",
    1554 => "110000100011",
    1555 => "110000100101",
    1556 => "110000100111",
    1557 => "110000101001",
    1558 => "110000101011",
    1559 => "110000101101",
    1560 => "110000101111",
    1561 => "110000110001",
    1562 => "110000110011",
    1563 => "110000110101",
    1564 => "110000110111",
    1565 => "110000111001",
    1566 => "110000111011",
    1567 => "110000111101",
    1568 => "110000111111",
    1569 => "110001000001",
    1570 => "110001000011",
    1571 => "110001000101",
    1572 => "110001000111",
    1573 => "110001001001",
    1574 => "110001001011",
    1575 => "110001001101",
    1576 => "110001001111",
    1577 => "110001010001",
    1578 => "110001010011",
    1579 => "110001010101",
    1580 => "110001010111",
    1581 => "110001011001",
    1582 => "110001011011",
    1583 => "110001011101",
    1584 => "110001011111",
    1585 => "110001100001",
    1586 => "110001100011",
    1587 => "110001100101",
    1588 => "110001100111",
    1589 => "110001101001",
    1590 => "110001101011",
    1591 => "110001101101",
    1592 => "110001101111",
    1593 => "110001110001",
    1594 => "110001110011",
    1595 => "110001110101",
    1596 => "110001110111",
    1597 => "110001111001",
    1598 => "110001111011",
    1599 => "110001111101",
    1600 => "110001111111",
    1601 => "110010000001",
    1602 => "110010000011",
    1603 => "110010000101",
    1604 => "110010000111",
    1605 => "110010001001",
    1606 => "110010001011",
    1607 => "110010001101",
    1608 => "110010001111",
    1609 => "110010010001",
    1610 => "110010010011",
    1611 => "110010010101",
    1612 => "110010010111",
    1613 => "110010011001",
    1614 => "110010011011",
    1615 => "110010011101",
    1616 => "110010011111",
    1617 => "110010100001",
    1618 => "110010100011",
    1619 => "110010100101",
    1620 => "110010100111",
    1621 => "110010101001",
    1622 => "110010101011",
    1623 => "110010101101",
    1624 => "110010101111",
    1625 => "110010110001",
    1626 => "110010110011",
    1627 => "110010110101",
    1628 => "110010110111",
    1629 => "110010111001",
    1630 => "110010111011",
    1631 => "110010111101",
    1632 => "110010111111",
    1633 => "110011000001",
    1634 => "110011000011",
    1635 => "110011000101",
    1636 => "110011000111",
    1637 => "110011001001",
    1638 => "110011001011",
    1639 => "110011001101",
    1640 => "110011001111",
    1641 => "110011010001",
    1642 => "110011010011",
    1643 => "110011010101",
    1644 => "110011010111",
    1645 => "110011011001",
    1646 => "110011011011",
    1647 => "110011011101",
    1648 => "110011011111",
    1649 => "110011100001",
    1650 => "110011100011",
    1651 => "110011100101",
    1652 => "110011100111",
    1653 => "110011101001",
    1654 => "110011101011",
    1655 => "110011101101",
    1656 => "110011101111",
    1657 => "110011110001",
    1658 => "110011110011",
    1659 => "110011110101",
    1660 => "110011110111",
    1661 => "110011111001",
    1662 => "110011111011",
    1663 => "110011111101",
    1664 => "110011111111",
    1665 => "110100000001",
    1666 => "110100000011",
    1667 => "110100000101",
    1668 => "110100000111",
    1669 => "110100001001",
    1670 => "110100001011",
    1671 => "110100001101",
    1672 => "110100001111",
    1673 => "110100010001",
    1674 => "110100010011",
    1675 => "110100010101",
    1676 => "110100010111",
    1677 => "110100011001",
    1678 => "110100011011",
    1679 => "110100011101",
    1680 => "110100011111",
    1681 => "110100100001",
    1682 => "110100100011",
    1683 => "110100100101",
    1684 => "110100100111",
    1685 => "110100101001",
    1686 => "110100101011",
    1687 => "110100101101",
    1688 => "110100101111",
    1689 => "110100110001",
    1690 => "110100110011",
    1691 => "110100110101",
    1692 => "110100110111",
    1693 => "110100111001",
    1694 => "110100111011",
    1695 => "110100111101",
    1696 => "110100111111",
    1697 => "110101000001",
    1698 => "110101000011",
    1699 => "110101000101",
    1700 => "110101000111",
    1701 => "110101001001",
    1702 => "110101001011",
    1703 => "110101001101",
    1704 => "110101001111",
    1705 => "110101010001",
    1706 => "110101010011",
    1707 => "110101010101",
    1708 => "110101010111",
    1709 => "110101011001",
    1710 => "110101011011",
    1711 => "110101011101",
    1712 => "110101011111",
    1713 => "110101100001",
    1714 => "110101100011",
    1715 => "110101100101",
    1716 => "110101100111",
    1717 => "110101101001",
    1718 => "110101101011",
    1719 => "110101101101",
    1720 => "110101101111",
    1721 => "110101110001",
    1722 => "110101110011",
    1723 => "110101110101",
    1724 => "110101110111",
    1725 => "110101111001",
    1726 => "110101111011",
    1727 => "110101111101",
    1728 => "110101111111",
    1729 => "110110000001",
    1730 => "110110000011",
    1731 => "110110000101",
    1732 => "110110000111",
    1733 => "110110001001",
    1734 => "110110001011",
    1735 => "110110001101",
    1736 => "110110001111",
    1737 => "110110010001",
    1738 => "110110010011",
    1739 => "110110010101",
    1740 => "110110010111",
    1741 => "110110011001",
    1742 => "110110011011",
    1743 => "110110011101",
    1744 => "110110011111",
    1745 => "110110100001",
    1746 => "110110100011",
    1747 => "110110100101",
    1748 => "110110100111",
    1749 => "110110101001",
    1750 => "110110101011",
    1751 => "110110101101",
    1752 => "110110101111",
    1753 => "110110110001",
    1754 => "110110110011",
    1755 => "110110110101",
    1756 => "110110110111",
    1757 => "110110111001",
    1758 => "110110111011",
    1759 => "110110111101",
    1760 => "110110111111",
    1761 => "110111000001",
    1762 => "110111000011",
    1763 => "110111000101",
    1764 => "110111000111",
    1765 => "110111001001",
    1766 => "110111001011",
    1767 => "110111001101",
    1768 => "110111001111",
    1769 => "110111010001",
    1770 => "110111010011",
    1771 => "110111010101",
    1772 => "110111010111",
    1773 => "110111011001",
    1774 => "110111011011",
    1775 => "110111011101",
    1776 => "110111011111",
    1777 => "110111100001",
    1778 => "110111100011",
    1779 => "110111100101",
    1780 => "110111100111",
    1781 => "110111101001",
    1782 => "110111101011",
    1783 => "110111101101",
    1784 => "110111101111",
    1785 => "110111110001",
    1786 => "110111110011",
    1787 => "110111110101",
    1788 => "110111110111",
    1789 => "110111111001",
    1790 => "110111111011",
    1791 => "110111111101",
    1792 => "110111111111",
    1793 => "111000000001",
    1794 => "111000000011",
    1795 => "111000000101",
    1796 => "111000000111",
    1797 => "111000001001",
    1798 => "111000001011",
    1799 => "111000001101",
    1800 => "111000001111",
    1801 => "111000010001",
    1802 => "111000010011",
    1803 => "111000010101",
    1804 => "111000010111",
    1805 => "111000011001",
    1806 => "111000011011",
    1807 => "111000011101",
    1808 => "111000011111",
    1809 => "111000100001",
    1810 => "111000100011",
    1811 => "111000100101",
    1812 => "111000100111",
    1813 => "111000101001",
    1814 => "111000101011",
    1815 => "111000101101",
    1816 => "111000101111",
    1817 => "111000110001",
    1818 => "111000110011",
    1819 => "111000110101",
    1820 => "111000110111",
    1821 => "111000111001",
    1822 => "111000111011",
    1823 => "111000111101",
    1824 => "111000111111",
    1825 => "111001000001",
    1826 => "111001000011",
    1827 => "111001000101",
    1828 => "111001000111",
    1829 => "111001001001",
    1830 => "111001001011",
    1831 => "111001001101",
    1832 => "111001001111",
    1833 => "111001010001",
    1834 => "111001010011",
    1835 => "111001010101",
    1836 => "111001010111",
    1837 => "111001011001",
    1838 => "111001011011",
    1839 => "111001011101",
    1840 => "111001011111",
    1841 => "111001100001",
    1842 => "111001100011",
    1843 => "111001100101",
    1844 => "111001100111",
    1845 => "111001101001",
    1846 => "111001101011",
    1847 => "111001101101",
    1848 => "111001101111",
    1849 => "111001110001",
    1850 => "111001110011",
    1851 => "111001110101",
    1852 => "111001110111",
    1853 => "111001111001",
    1854 => "111001111011",
    1855 => "111001111101",
    1856 => "111001111111",
    1857 => "111010000001",
    1858 => "111010000011",
    1859 => "111010000101",
    1860 => "111010000111",
    1861 => "111010001001",
    1862 => "111010001011",
    1863 => "111010001101",
    1864 => "111010001111",
    1865 => "111010010001",
    1866 => "111010010011",
    1867 => "111010010101",
    1868 => "111010010111",
    1869 => "111010011001",
    1870 => "111010011011",
    1871 => "111010011101",
    1872 => "111010011111",
    1873 => "111010100001",
    1874 => "111010100011",
    1875 => "111010100101",
    1876 => "111010100111",
    1877 => "111010101001",
    1878 => "111010101011",
    1879 => "111010101101",
    1880 => "111010101111",
    1881 => "111010110001",
    1882 => "111010110011",
    1883 => "111010110101",
    1884 => "111010110111",
    1885 => "111010111001",
    1886 => "111010111011",
    1887 => "111010111101",
    1888 => "111010111111",
    1889 => "111011000001",
    1890 => "111011000011",
    1891 => "111011000101",
    1892 => "111011000111",
    1893 => "111011001001",
    1894 => "111011001011",
    1895 => "111011001101",
    1896 => "111011001111",
    1897 => "111011010001",
    1898 => "111011010011",
    1899 => "111011010101",
    1900 => "111011010111",
    1901 => "111011011001",
    1902 => "111011011011",
    1903 => "111011011101",
    1904 => "111011011111",
    1905 => "111011100001",
    1906 => "111011100011",
    1907 => "111011100101",
    1908 => "111011100111",
    1909 => "111011101001",
    1910 => "111011101011",
    1911 => "111011101101",
    1912 => "111011101111",
    1913 => "111011110001",
    1914 => "111011110011",
    1915 => "111011110101",
    1916 => "111011110111",
    1917 => "111011111001",
    1918 => "111011111011",
    1919 => "111011111101",
    1920 => "111011111111",
    1921 => "111100000001",
    1922 => "111100000011",
    1923 => "111100000101",
    1924 => "111100000111",
    1925 => "111100001001",
    1926 => "111100001011",
    1927 => "111100001101",
    1928 => "111100001111",
    1929 => "111100010001",
    1930 => "111100010011",
    1931 => "111100010101",
    1932 => "111100010111",
    1933 => "111100011001",
    1934 => "111100011011",
    1935 => "111100011101",
    1936 => "111100011111",
    1937 => "111100100001",
    1938 => "111100100011",
    1939 => "111100100101",
    1940 => "111100100111",
    1941 => "111100101001",
    1942 => "111100101011",
    1943 => "111100101101",
    1944 => "111100101111",
    1945 => "111100110001",
    1946 => "111100110011",
    1947 => "111100110101",
    1948 => "111100110111",
    1949 => "111100111001",
    1950 => "111100111011",
    1951 => "111100111101",
    1952 => "111100111111",
    1953 => "111101000001",
    1954 => "111101000011",
    1955 => "111101000101",
    1956 => "111101000111",
    1957 => "111101001001",
    1958 => "111101001011",
    1959 => "111101001101",
    1960 => "111101001111",
    1961 => "111101010001",
    1962 => "111101010011",
    1963 => "111101010101",
    1964 => "111101010111",
    1965 => "111101011001",
    1966 => "111101011011",
    1967 => "111101011101",
    1968 => "111101011111",
    1969 => "111101100001",
    1970 => "111101100011",
    1971 => "111101100101",
    1972 => "111101100111",
    1973 => "111101101001",
    1974 => "111101101011",
    1975 => "111101101101",
    1976 => "111101101111",
    1977 => "111101110001",
    1978 => "111101110011",
    1979 => "111101110101",
    1980 => "111101110111",
    1981 => "111101111001",
    1982 => "111101111011",
    1983 => "111101111101",
    1984 => "111101111111",
    1985 => "111110000001",
    1986 => "111110000011",
    1987 => "111110000101",
    1988 => "111110000111",
    1989 => "111110001001",
    1990 => "111110001011",
    1991 => "111110001101",
    1992 => "111110001111",
    1993 => "111110010001",
    1994 => "111110010011",
    1995 => "111110010101",
    1996 => "111110010111",
    1997 => "111110011001",
    1998 => "111110011011",
    1999 => "111110011101",
    2000 => "111110011111",
    2001 => "111110100001",
    2002 => "111110100011",
    2003 => "111110100101",
    2004 => "111110100111",
    2005 => "111110101001",
    2006 => "111110101011",
    2007 => "111110101101",
    2008 => "111110101111",
    2009 => "111110110001",
    2010 => "111110110011",
    2011 => "111110110101",
    2012 => "111110110111",
    2013 => "111110111001",
    2014 => "111110111011",
    2015 => "111110111101",
    2016 => "111110111111",
    2017 => "111111000001",
    2018 => "111111000011",
    2019 => "111111000101",
    2020 => "111111000111",
    2021 => "111111001001",
    2022 => "111111001011",
    2023 => "111111001101",
    2024 => "111111001111",
    2025 => "111111010001",
    2026 => "111111010011",
    2027 => "111111010101",
    2028 => "111111010111",
    2029 => "111111011001",
    2030 => "111111011011",
    2031 => "111111011101",
    2032 => "111111011111",
    2033 => "111111100001",
    2034 => "111111100011",
    2035 => "111111100101",
    2036 => "111111100111",
    2037 => "111111101001",
    2038 => "111111101011",
    2039 => "111111101101",
    2040 => "111111101111",
    2041 => "111111110001",
    2042 => "111111110011",
    2043 => "111111110101",
    2044 => "111111110111",
    2045 => "111111111001",
    2046 => "111111111011",
    2047 => "111111111101",
    2048 => "111111111111",
    2049 => "111111111101",
    2050 => "111111111011",
    2051 => "111111111001",
    2052 => "111111110111",
    2053 => "111111110101",
    2054 => "111111110011",
    2055 => "111111110001",
    2056 => "111111101111",
    2057 => "111111101101",
    2058 => "111111101011",
    2059 => "111111101001",
    2060 => "111111100111",
    2061 => "111111100101",
    2062 => "111111100011",
    2063 => "111111100001",
    2064 => "111111011111",
    2065 => "111111011101",
    2066 => "111111011011",
    2067 => "111111011001",
    2068 => "111111010111",
    2069 => "111111010101",
    2070 => "111111010011",
    2071 => "111111010001",
    2072 => "111111001111",
    2073 => "111111001101",
    2074 => "111111001011",
    2075 => "111111001001",
    2076 => "111111000111",
    2077 => "111111000101",
    2078 => "111111000011",
    2079 => "111111000001",
    2080 => "111110111111",
    2081 => "111110111101",
    2082 => "111110111011",
    2083 => "111110111001",
    2084 => "111110110111",
    2085 => "111110110101",
    2086 => "111110110011",
    2087 => "111110110001",
    2088 => "111110101111",
    2089 => "111110101101",
    2090 => "111110101011",
    2091 => "111110101001",
    2092 => "111110100111",
    2093 => "111110100101",
    2094 => "111110100011",
    2095 => "111110100001",
    2096 => "111110011111",
    2097 => "111110011101",
    2098 => "111110011011",
    2099 => "111110011001",
    2100 => "111110010111",
    2101 => "111110010101",
    2102 => "111110010011",
    2103 => "111110010001",
    2104 => "111110001111",
    2105 => "111110001101",
    2106 => "111110001011",
    2107 => "111110001001",
    2108 => "111110000111",
    2109 => "111110000101",
    2110 => "111110000011",
    2111 => "111110000001",
    2112 => "111101111111",
    2113 => "111101111101",
    2114 => "111101111011",
    2115 => "111101111001",
    2116 => "111101110111",
    2117 => "111101110101",
    2118 => "111101110011",
    2119 => "111101110001",
    2120 => "111101101111",
    2121 => "111101101101",
    2122 => "111101101011",
    2123 => "111101101001",
    2124 => "111101100111",
    2125 => "111101100101",
    2126 => "111101100011",
    2127 => "111101100001",
    2128 => "111101011111",
    2129 => "111101011101",
    2130 => "111101011011",
    2131 => "111101011001",
    2132 => "111101010111",
    2133 => "111101010101",
    2134 => "111101010011",
    2135 => "111101010001",
    2136 => "111101001111",
    2137 => "111101001101",
    2138 => "111101001011",
    2139 => "111101001001",
    2140 => "111101000111",
    2141 => "111101000101",
    2142 => "111101000011",
    2143 => "111101000001",
    2144 => "111100111111",
    2145 => "111100111101",
    2146 => "111100111011",
    2147 => "111100111001",
    2148 => "111100110111",
    2149 => "111100110101",
    2150 => "111100110011",
    2151 => "111100110001",
    2152 => "111100101111",
    2153 => "111100101101",
    2154 => "111100101011",
    2155 => "111100101001",
    2156 => "111100100111",
    2157 => "111100100101",
    2158 => "111100100011",
    2159 => "111100100001",
    2160 => "111100011111",
    2161 => "111100011101",
    2162 => "111100011011",
    2163 => "111100011001",
    2164 => "111100010111",
    2165 => "111100010101",
    2166 => "111100010011",
    2167 => "111100010001",
    2168 => "111100001111",
    2169 => "111100001101",
    2170 => "111100001011",
    2171 => "111100001001",
    2172 => "111100000111",
    2173 => "111100000101",
    2174 => "111100000011",
    2175 => "111100000001",
    2176 => "111011111111",
    2177 => "111011111101",
    2178 => "111011111011",
    2179 => "111011111001",
    2180 => "111011110111",
    2181 => "111011110101",
    2182 => "111011110011",
    2183 => "111011110001",
    2184 => "111011101111",
    2185 => "111011101101",
    2186 => "111011101011",
    2187 => "111011101001",
    2188 => "111011100111",
    2189 => "111011100101",
    2190 => "111011100011",
    2191 => "111011100001",
    2192 => "111011011111",
    2193 => "111011011101",
    2194 => "111011011011",
    2195 => "111011011001",
    2196 => "111011010111",
    2197 => "111011010101",
    2198 => "111011010011",
    2199 => "111011010001",
    2200 => "111011001111",
    2201 => "111011001101",
    2202 => "111011001011",
    2203 => "111011001001",
    2204 => "111011000111",
    2205 => "111011000101",
    2206 => "111011000011",
    2207 => "111011000001",
    2208 => "111010111111",
    2209 => "111010111101",
    2210 => "111010111011",
    2211 => "111010111001",
    2212 => "111010110111",
    2213 => "111010110101",
    2214 => "111010110011",
    2215 => "111010110001",
    2216 => "111010101111",
    2217 => "111010101101",
    2218 => "111010101011",
    2219 => "111010101001",
    2220 => "111010100111",
    2221 => "111010100101",
    2222 => "111010100011",
    2223 => "111010100001",
    2224 => "111010011111",
    2225 => "111010011101",
    2226 => "111010011011",
    2227 => "111010011001",
    2228 => "111010010111",
    2229 => "111010010101",
    2230 => "111010010011",
    2231 => "111010010001",
    2232 => "111010001111",
    2233 => "111010001101",
    2234 => "111010001011",
    2235 => "111010001001",
    2236 => "111010000111",
    2237 => "111010000101",
    2238 => "111010000011",
    2239 => "111010000001",
    2240 => "111001111111",
    2241 => "111001111101",
    2242 => "111001111011",
    2243 => "111001111001",
    2244 => "111001110111",
    2245 => "111001110101",
    2246 => "111001110011",
    2247 => "111001110001",
    2248 => "111001101111",
    2249 => "111001101101",
    2250 => "111001101011",
    2251 => "111001101001",
    2252 => "111001100111",
    2253 => "111001100101",
    2254 => "111001100011",
    2255 => "111001100001",
    2256 => "111001011111",
    2257 => "111001011101",
    2258 => "111001011011",
    2259 => "111001011001",
    2260 => "111001010111",
    2261 => "111001010101",
    2262 => "111001010011",
    2263 => "111001010001",
    2264 => "111001001111",
    2265 => "111001001101",
    2266 => "111001001011",
    2267 => "111001001001",
    2268 => "111001000111",
    2269 => "111001000101",
    2270 => "111001000011",
    2271 => "111001000001",
    2272 => "111000111111",
    2273 => "111000111101",
    2274 => "111000111011",
    2275 => "111000111001",
    2276 => "111000110111",
    2277 => "111000110101",
    2278 => "111000110011",
    2279 => "111000110001",
    2280 => "111000101111",
    2281 => "111000101101",
    2282 => "111000101011",
    2283 => "111000101001",
    2284 => "111000100111",
    2285 => "111000100101",
    2286 => "111000100011",
    2287 => "111000100001",
    2288 => "111000011111",
    2289 => "111000011101",
    2290 => "111000011011",
    2291 => "111000011001",
    2292 => "111000010111",
    2293 => "111000010101",
    2294 => "111000010011",
    2295 => "111000010001",
    2296 => "111000001111",
    2297 => "111000001101",
    2298 => "111000001011",
    2299 => "111000001001",
    2300 => "111000000111",
    2301 => "111000000101",
    2302 => "111000000011",
    2303 => "111000000001",
    2304 => "110111111111",
    2305 => "110111111101",
    2306 => "110111111011",
    2307 => "110111111001",
    2308 => "110111110111",
    2309 => "110111110101",
    2310 => "110111110011",
    2311 => "110111110001",
    2312 => "110111101111",
    2313 => "110111101101",
    2314 => "110111101011",
    2315 => "110111101001",
    2316 => "110111100111",
    2317 => "110111100101",
    2318 => "110111100011",
    2319 => "110111100001",
    2320 => "110111011111",
    2321 => "110111011101",
    2322 => "110111011011",
    2323 => "110111011001",
    2324 => "110111010111",
    2325 => "110111010101",
    2326 => "110111010011",
    2327 => "110111010001",
    2328 => "110111001111",
    2329 => "110111001101",
    2330 => "110111001011",
    2331 => "110111001001",
    2332 => "110111000111",
    2333 => "110111000101",
    2334 => "110111000011",
    2335 => "110111000001",
    2336 => "110110111111",
    2337 => "110110111101",
    2338 => "110110111011",
    2339 => "110110111001",
    2340 => "110110110111",
    2341 => "110110110101",
    2342 => "110110110011",
    2343 => "110110110001",
    2344 => "110110101111",
    2345 => "110110101101",
    2346 => "110110101011",
    2347 => "110110101001",
    2348 => "110110100111",
    2349 => "110110100101",
    2350 => "110110100011",
    2351 => "110110100001",
    2352 => "110110011111",
    2353 => "110110011101",
    2354 => "110110011011",
    2355 => "110110011001",
    2356 => "110110010111",
    2357 => "110110010101",
    2358 => "110110010011",
    2359 => "110110010001",
    2360 => "110110001111",
    2361 => "110110001101",
    2362 => "110110001011",
    2363 => "110110001001",
    2364 => "110110000111",
    2365 => "110110000101",
    2366 => "110110000011",
    2367 => "110110000001",
    2368 => "110101111111",
    2369 => "110101111101",
    2370 => "110101111011",
    2371 => "110101111001",
    2372 => "110101110111",
    2373 => "110101110101",
    2374 => "110101110011",
    2375 => "110101110001",
    2376 => "110101101111",
    2377 => "110101101101",
    2378 => "110101101011",
    2379 => "110101101001",
    2380 => "110101100111",
    2381 => "110101100101",
    2382 => "110101100011",
    2383 => "110101100001",
    2384 => "110101011111",
    2385 => "110101011101",
    2386 => "110101011011",
    2387 => "110101011001",
    2388 => "110101010111",
    2389 => "110101010101",
    2390 => "110101010011",
    2391 => "110101010001",
    2392 => "110101001111",
    2393 => "110101001101",
    2394 => "110101001011",
    2395 => "110101001001",
    2396 => "110101000111",
    2397 => "110101000101",
    2398 => "110101000011",
    2399 => "110101000001",
    2400 => "110100111111",
    2401 => "110100111101",
    2402 => "110100111011",
    2403 => "110100111001",
    2404 => "110100110111",
    2405 => "110100110101",
    2406 => "110100110011",
    2407 => "110100110001",
    2408 => "110100101111",
    2409 => "110100101101",
    2410 => "110100101011",
    2411 => "110100101001",
    2412 => "110100100111",
    2413 => "110100100101",
    2414 => "110100100011",
    2415 => "110100100001",
    2416 => "110100011111",
    2417 => "110100011101",
    2418 => "110100011011",
    2419 => "110100011001",
    2420 => "110100010111",
    2421 => "110100010101",
    2422 => "110100010011",
    2423 => "110100010001",
    2424 => "110100001111",
    2425 => "110100001101",
    2426 => "110100001011",
    2427 => "110100001001",
    2428 => "110100000111",
    2429 => "110100000101",
    2430 => "110100000011",
    2431 => "110100000001",
    2432 => "110011111111",
    2433 => "110011111101",
    2434 => "110011111011",
    2435 => "110011111001",
    2436 => "110011110111",
    2437 => "110011110101",
    2438 => "110011110011",
    2439 => "110011110001",
    2440 => "110011101111",
    2441 => "110011101101",
    2442 => "110011101011",
    2443 => "110011101001",
    2444 => "110011100111",
    2445 => "110011100101",
    2446 => "110011100011",
    2447 => "110011100001",
    2448 => "110011011111",
    2449 => "110011011101",
    2450 => "110011011011",
    2451 => "110011011001",
    2452 => "110011010111",
    2453 => "110011010101",
    2454 => "110011010011",
    2455 => "110011010001",
    2456 => "110011001111",
    2457 => "110011001101",
    2458 => "110011001011",
    2459 => "110011001001",
    2460 => "110011000111",
    2461 => "110011000101",
    2462 => "110011000011",
    2463 => "110011000001",
    2464 => "110010111111",
    2465 => "110010111101",
    2466 => "110010111011",
    2467 => "110010111001",
    2468 => "110010110111",
    2469 => "110010110101",
    2470 => "110010110011",
    2471 => "110010110001",
    2472 => "110010101111",
    2473 => "110010101101",
    2474 => "110010101011",
    2475 => "110010101001",
    2476 => "110010100111",
    2477 => "110010100101",
    2478 => "110010100011",
    2479 => "110010100001",
    2480 => "110010011111",
    2481 => "110010011101",
    2482 => "110010011011",
    2483 => "110010011001",
    2484 => "110010010111",
    2485 => "110010010101",
    2486 => "110010010011",
    2487 => "110010010001",
    2488 => "110010001111",
    2489 => "110010001101",
    2490 => "110010001011",
    2491 => "110010001001",
    2492 => "110010000111",
    2493 => "110010000101",
    2494 => "110010000011",
    2495 => "110010000001",
    2496 => "110001111111",
    2497 => "110001111101",
    2498 => "110001111011",
    2499 => "110001111001",
    2500 => "110001110111",
    2501 => "110001110101",
    2502 => "110001110011",
    2503 => "110001110001",
    2504 => "110001101111",
    2505 => "110001101101",
    2506 => "110001101011",
    2507 => "110001101001",
    2508 => "110001100111",
    2509 => "110001100101",
    2510 => "110001100011",
    2511 => "110001100001",
    2512 => "110001011111",
    2513 => "110001011101",
    2514 => "110001011011",
    2515 => "110001011001",
    2516 => "110001010111",
    2517 => "110001010101",
    2518 => "110001010011",
    2519 => "110001010001",
    2520 => "110001001111",
    2521 => "110001001101",
    2522 => "110001001011",
    2523 => "110001001001",
    2524 => "110001000111",
    2525 => "110001000101",
    2526 => "110001000011",
    2527 => "110001000001",
    2528 => "110000111111",
    2529 => "110000111101",
    2530 => "110000111011",
    2531 => "110000111001",
    2532 => "110000110111",
    2533 => "110000110101",
    2534 => "110000110011",
    2535 => "110000110001",
    2536 => "110000101111",
    2537 => "110000101101",
    2538 => "110000101011",
    2539 => "110000101001",
    2540 => "110000100111",
    2541 => "110000100101",
    2542 => "110000100011",
    2543 => "110000100001",
    2544 => "110000011111",
    2545 => "110000011101",
    2546 => "110000011011",
    2547 => "110000011001",
    2548 => "110000010111",
    2549 => "110000010101",
    2550 => "110000010011",
    2551 => "110000010001",
    2552 => "110000001111",
    2553 => "110000001101",
    2554 => "110000001011",
    2555 => "110000001001",
    2556 => "110000000111",
    2557 => "110000000101",
    2558 => "110000000011",
    2559 => "110000000001",
    2560 => "101111111111",
    2561 => "101111111101",
    2562 => "101111111011",
    2563 => "101111111001",
    2564 => "101111110111",
    2565 => "101111110101",
    2566 => "101111110011",
    2567 => "101111110001",
    2568 => "101111101111",
    2569 => "101111101101",
    2570 => "101111101011",
    2571 => "101111101001",
    2572 => "101111100111",
    2573 => "101111100101",
    2574 => "101111100011",
    2575 => "101111100001",
    2576 => "101111011111",
    2577 => "101111011101",
    2578 => "101111011011",
    2579 => "101111011001",
    2580 => "101111010111",
    2581 => "101111010101",
    2582 => "101111010011",
    2583 => "101111010001",
    2584 => "101111001111",
    2585 => "101111001101",
    2586 => "101111001011",
    2587 => "101111001001",
    2588 => "101111000111",
    2589 => "101111000101",
    2590 => "101111000011",
    2591 => "101111000001",
    2592 => "101110111111",
    2593 => "101110111101",
    2594 => "101110111011",
    2595 => "101110111001",
    2596 => "101110110111",
    2597 => "101110110101",
    2598 => "101110110011",
    2599 => "101110110001",
    2600 => "101110101111",
    2601 => "101110101101",
    2602 => "101110101011",
    2603 => "101110101001",
    2604 => "101110100111",
    2605 => "101110100101",
    2606 => "101110100011",
    2607 => "101110100001",
    2608 => "101110011111",
    2609 => "101110011101",
    2610 => "101110011011",
    2611 => "101110011001",
    2612 => "101110010111",
    2613 => "101110010101",
    2614 => "101110010011",
    2615 => "101110010001",
    2616 => "101110001111",
    2617 => "101110001101",
    2618 => "101110001011",
    2619 => "101110001001",
    2620 => "101110000111",
    2621 => "101110000101",
    2622 => "101110000011",
    2623 => "101110000001",
    2624 => "101101111111",
    2625 => "101101111101",
    2626 => "101101111011",
    2627 => "101101111001",
    2628 => "101101110111",
    2629 => "101101110101",
    2630 => "101101110011",
    2631 => "101101110001",
    2632 => "101101101111",
    2633 => "101101101101",
    2634 => "101101101011",
    2635 => "101101101001",
    2636 => "101101100111",
    2637 => "101101100101",
    2638 => "101101100011",
    2639 => "101101100001",
    2640 => "101101011111",
    2641 => "101101011101",
    2642 => "101101011011",
    2643 => "101101011001",
    2644 => "101101010111",
    2645 => "101101010101",
    2646 => "101101010011",
    2647 => "101101010001",
    2648 => "101101001111",
    2649 => "101101001101",
    2650 => "101101001011",
    2651 => "101101001001",
    2652 => "101101000111",
    2653 => "101101000101",
    2654 => "101101000011",
    2655 => "101101000001",
    2656 => "101100111111",
    2657 => "101100111101",
    2658 => "101100111011",
    2659 => "101100111001",
    2660 => "101100110111",
    2661 => "101100110101",
    2662 => "101100110011",
    2663 => "101100110001",
    2664 => "101100101111",
    2665 => "101100101101",
    2666 => "101100101011",
    2667 => "101100101001",
    2668 => "101100100111",
    2669 => "101100100101",
    2670 => "101100100011",
    2671 => "101100100001",
    2672 => "101100011111",
    2673 => "101100011101",
    2674 => "101100011011",
    2675 => "101100011001",
    2676 => "101100010111",
    2677 => "101100010101",
    2678 => "101100010011",
    2679 => "101100010001",
    2680 => "101100001111",
    2681 => "101100001101",
    2682 => "101100001011",
    2683 => "101100001001",
    2684 => "101100000111",
    2685 => "101100000101",
    2686 => "101100000011",
    2687 => "101100000001",
    2688 => "101011111111",
    2689 => "101011111101",
    2690 => "101011111011",
    2691 => "101011111001",
    2692 => "101011110111",
    2693 => "101011110101",
    2694 => "101011110011",
    2695 => "101011110001",
    2696 => "101011101111",
    2697 => "101011101101",
    2698 => "101011101011",
    2699 => "101011101001",
    2700 => "101011100111",
    2701 => "101011100101",
    2702 => "101011100011",
    2703 => "101011100001",
    2704 => "101011011111",
    2705 => "101011011101",
    2706 => "101011011011",
    2707 => "101011011001",
    2708 => "101011010111",
    2709 => "101011010101",
    2710 => "101011010011",
    2711 => "101011010001",
    2712 => "101011001111",
    2713 => "101011001101",
    2714 => "101011001011",
    2715 => "101011001001",
    2716 => "101011000111",
    2717 => "101011000101",
    2718 => "101011000011",
    2719 => "101011000001",
    2720 => "101010111111",
    2721 => "101010111101",
    2722 => "101010111011",
    2723 => "101010111001",
    2724 => "101010110111",
    2725 => "101010110101",
    2726 => "101010110011",
    2727 => "101010110001",
    2728 => "101010101111",
    2729 => "101010101101",
    2730 => "101010101011",
    2731 => "101010101001",
    2732 => "101010100111",
    2733 => "101010100101",
    2734 => "101010100011",
    2735 => "101010100001",
    2736 => "101010011111",
    2737 => "101010011101",
    2738 => "101010011011",
    2739 => "101010011001",
    2740 => "101010010111",
    2741 => "101010010101",
    2742 => "101010010011",
    2743 => "101010010001",
    2744 => "101010001111",
    2745 => "101010001101",
    2746 => "101010001011",
    2747 => "101010001001",
    2748 => "101010000111",
    2749 => "101010000101",
    2750 => "101010000011",
    2751 => "101010000001",
    2752 => "101001111111",
    2753 => "101001111101",
    2754 => "101001111011",
    2755 => "101001111001",
    2756 => "101001110111",
    2757 => "101001110101",
    2758 => "101001110011",
    2759 => "101001110001",
    2760 => "101001101111",
    2761 => "101001101101",
    2762 => "101001101011",
    2763 => "101001101001",
    2764 => "101001100111",
    2765 => "101001100101",
    2766 => "101001100011",
    2767 => "101001100001",
    2768 => "101001011111",
    2769 => "101001011101",
    2770 => "101001011011",
    2771 => "101001011001",
    2772 => "101001010111",
    2773 => "101001010101",
    2774 => "101001010011",
    2775 => "101001010001",
    2776 => "101001001111",
    2777 => "101001001101",
    2778 => "101001001011",
    2779 => "101001001001",
    2780 => "101001000111",
    2781 => "101001000101",
    2782 => "101001000011",
    2783 => "101001000001",
    2784 => "101000111111",
    2785 => "101000111101",
    2786 => "101000111011",
    2787 => "101000111001",
    2788 => "101000110111",
    2789 => "101000110101",
    2790 => "101000110011",
    2791 => "101000110001",
    2792 => "101000101111",
    2793 => "101000101101",
    2794 => "101000101011",
    2795 => "101000101001",
    2796 => "101000100111",
    2797 => "101000100101",
    2798 => "101000100011",
    2799 => "101000100001",
    2800 => "101000011111",
    2801 => "101000011101",
    2802 => "101000011011",
    2803 => "101000011001",
    2804 => "101000010111",
    2805 => "101000010101",
    2806 => "101000010011",
    2807 => "101000010001",
    2808 => "101000001111",
    2809 => "101000001101",
    2810 => "101000001011",
    2811 => "101000001001",
    2812 => "101000000111",
    2813 => "101000000101",
    2814 => "101000000011",
    2815 => "101000000001",
    2816 => "100111111111",
    2817 => "100111111101",
    2818 => "100111111011",
    2819 => "100111111001",
    2820 => "100111110111",
    2821 => "100111110101",
    2822 => "100111110011",
    2823 => "100111110001",
    2824 => "100111101111",
    2825 => "100111101101",
    2826 => "100111101011",
    2827 => "100111101001",
    2828 => "100111100111",
    2829 => "100111100101",
    2830 => "100111100011",
    2831 => "100111100001",
    2832 => "100111011111",
    2833 => "100111011101",
    2834 => "100111011011",
    2835 => "100111011001",
    2836 => "100111010111",
    2837 => "100111010101",
    2838 => "100111010011",
    2839 => "100111010001",
    2840 => "100111001111",
    2841 => "100111001101",
    2842 => "100111001011",
    2843 => "100111001001",
    2844 => "100111000111",
    2845 => "100111000101",
    2846 => "100111000100",
    2847 => "100111000010",
    2848 => "100111000000",
    2849 => "100110111110",
    2850 => "100110111100",
    2851 => "100110111010",
    2852 => "100110111000",
    2853 => "100110110110",
    2854 => "100110110100",
    2855 => "100110110010",
    2856 => "100110110000",
    2857 => "100110101110",
    2858 => "100110101100",
    2859 => "100110101010",
    2860 => "100110101000",
    2861 => "100110100110",
    2862 => "100110100100",
    2863 => "100110100010",
    2864 => "100110100000",
    2865 => "100110011110",
    2866 => "100110011100",
    2867 => "100110011010",
    2868 => "100110011000",
    2869 => "100110010110",
    2870 => "100110010100",
    2871 => "100110010010",
    2872 => "100110010000",
    2873 => "100110001110",
    2874 => "100110001100",
    2875 => "100110001010",
    2876 => "100110001000",
    2877 => "100110000110",
    2878 => "100110000100",
    2879 => "100110000010",
    2880 => "100110000000",
    2881 => "100101111110",
    2882 => "100101111100",
    2883 => "100101111010",
    2884 => "100101111000",
    2885 => "100101110110",
    2886 => "100101110100",
    2887 => "100101110010",
    2888 => "100101110000",
    2889 => "100101101110",
    2890 => "100101101100",
    2891 => "100101101010",
    2892 => "100101101000",
    2893 => "100101100110",
    2894 => "100101100100",
    2895 => "100101100010",
    2896 => "100101100000",
    2897 => "100101011110",
    2898 => "100101011100",
    2899 => "100101011010",
    2900 => "100101011000",
    2901 => "100101010110",
    2902 => "100101010100",
    2903 => "100101010010",
    2904 => "100101010000",
    2905 => "100101001110",
    2906 => "100101001100",
    2907 => "100101001010",
    2908 => "100101001000",
    2909 => "100101000110",
    2910 => "100101000100",
    2911 => "100101000010",
    2912 => "100101000000",
    2913 => "100100111110",
    2914 => "100100111100",
    2915 => "100100111010",
    2916 => "100100111000",
    2917 => "100100110110",
    2918 => "100100110100",
    2919 => "100100110010",
    2920 => "100100110000",
    2921 => "100100101110",
    2922 => "100100101100",
    2923 => "100100101010",
    2924 => "100100101000",
    2925 => "100100100110",
    2926 => "100100100100",
    2927 => "100100100010",
    2928 => "100100100000",
    2929 => "100100011110",
    2930 => "100100011100",
    2931 => "100100011010",
    2932 => "100100011000",
    2933 => "100100010110",
    2934 => "100100010100",
    2935 => "100100010010",
    2936 => "100100010000",
    2937 => "100100001110",
    2938 => "100100001100",
    2939 => "100100001010",
    2940 => "100100001000",
    2941 => "100100000110",
    2942 => "100100000100",
    2943 => "100100000010",
    2944 => "100100000000",
    2945 => "100011111110",
    2946 => "100011111100",
    2947 => "100011111010",
    2948 => "100011111000",
    2949 => "100011110110",
    2950 => "100011110100",
    2951 => "100011110010",
    2952 => "100011110000",
    2953 => "100011101110",
    2954 => "100011101100",
    2955 => "100011101010",
    2956 => "100011101000",
    2957 => "100011100110",
    2958 => "100011100100",
    2959 => "100011100010",
    2960 => "100011100000",
    2961 => "100011011110",
    2962 => "100011011100",
    2963 => "100011011010",
    2964 => "100011011000",
    2965 => "100011010110",
    2966 => "100011010100",
    2967 => "100011010010",
    2968 => "100011010000",
    2969 => "100011001110",
    2970 => "100011001100",
    2971 => "100011001010",
    2972 => "100011001000",
    2973 => "100011000110",
    2974 => "100011000100",
    2975 => "100011000010",
    2976 => "100011000000",
    2977 => "100010111110",
    2978 => "100010111100",
    2979 => "100010111010",
    2980 => "100010111000",
    2981 => "100010110110",
    2982 => "100010110100",
    2983 => "100010110010",
    2984 => "100010110000",
    2985 => "100010101110",
    2986 => "100010101100",
    2987 => "100010101010",
    2988 => "100010101000",
    2989 => "100010100110",
    2990 => "100010100100",
    2991 => "100010100010",
    2992 => "100010100000",
    2993 => "100010011110",
    2994 => "100010011100",
    2995 => "100010011010",
    2996 => "100010011000",
    2997 => "100010010110",
    2998 => "100010010100",
    2999 => "100010010010",
    3000 => "100010010000",
    3001 => "100010001110",
    3002 => "100010001100",
    3003 => "100010001010",
    3004 => "100010001000",
    3005 => "100010000110",
    3006 => "100010000100",
    3007 => "100010000010",
    3008 => "100010000000",
    3009 => "100001111110",
    3010 => "100001111100",
    3011 => "100001111010",
    3012 => "100001111000",
    3013 => "100001110110",
    3014 => "100001110100",
    3015 => "100001110010",
    3016 => "100001110000",
    3017 => "100001101110",
    3018 => "100001101100",
    3019 => "100001101010",
    3020 => "100001101000",
    3021 => "100001100110",
    3022 => "100001100100",
    3023 => "100001100010",
    3024 => "100001100000",
    3025 => "100001011110",
    3026 => "100001011100",
    3027 => "100001011010",
    3028 => "100001011000",
    3029 => "100001010110",
    3030 => "100001010100",
    3031 => "100001010010",
    3032 => "100001010000",
    3033 => "100001001110",
    3034 => "100001001100",
    3035 => "100001001010",
    3036 => "100001001000",
    3037 => "100001000110",
    3038 => "100001000100",
    3039 => "100001000010",
    3040 => "100001000000",
    3041 => "100000111110",
    3042 => "100000111100",
    3043 => "100000111010",
    3044 => "100000111000",
    3045 => "100000110110",
    3046 => "100000110100",
    3047 => "100000110010",
    3048 => "100000110000",
    3049 => "100000101110",
    3050 => "100000101100",
    3051 => "100000101010",
    3052 => "100000101000",
    3053 => "100000100110",
    3054 => "100000100100",
    3055 => "100000100010",
    3056 => "100000100000",
    3057 => "100000011110",
    3058 => "100000011100",
    3059 => "100000011010",
    3060 => "100000011000",
    3061 => "100000010110",
    3062 => "100000010100",
    3063 => "100000010010",
    3064 => "100000010000",
    3065 => "100000001110",
    3066 => "100000001100",
    3067 => "100000001010",
    3068 => "100000001000",
    3069 => "100000000110",
    3070 => "100000000100",
    3071 => "100000000010",
    3072 => "100000000000",
    3073 => "011111111110",
    3074 => "011111111100",
    3075 => "011111111010",
    3076 => "011111111000",
    3077 => "011111110110",
    3078 => "011111110100",
    3079 => "011111110010",
    3080 => "011111110000",
    3081 => "011111101110",
    3082 => "011111101100",
    3083 => "011111101010",
    3084 => "011111101000",
    3085 => "011111100110",
    3086 => "011111100100",
    3087 => "011111100010",
    3088 => "011111100000",
    3089 => "011111011110",
    3090 => "011111011100",
    3091 => "011111011010",
    3092 => "011111011000",
    3093 => "011111010110",
    3094 => "011111010100",
    3095 => "011111010010",
    3096 => "011111010000",
    3097 => "011111001110",
    3098 => "011111001100",
    3099 => "011111001010",
    3100 => "011111001000",
    3101 => "011111000110",
    3102 => "011111000100",
    3103 => "011111000010",
    3104 => "011111000000",
    3105 => "011110111110",
    3106 => "011110111100",
    3107 => "011110111010",
    3108 => "011110111000",
    3109 => "011110110110",
    3110 => "011110110100",
    3111 => "011110110010",
    3112 => "011110110000",
    3113 => "011110101110",
    3114 => "011110101100",
    3115 => "011110101010",
    3116 => "011110101000",
    3117 => "011110100110",
    3118 => "011110100100",
    3119 => "011110100010",
    3120 => "011110100000",
    3121 => "011110011110",
    3122 => "011110011100",
    3123 => "011110011010",
    3124 => "011110011000",
    3125 => "011110010110",
    3126 => "011110010100",
    3127 => "011110010010",
    3128 => "011110010000",
    3129 => "011110001110",
    3130 => "011110001100",
    3131 => "011110001010",
    3132 => "011110001000",
    3133 => "011110000110",
    3134 => "011110000100",
    3135 => "011110000010",
    3136 => "011110000000",
    3137 => "011101111110",
    3138 => "011101111100",
    3139 => "011101111010",
    3140 => "011101111000",
    3141 => "011101110110",
    3142 => "011101110100",
    3143 => "011101110010",
    3144 => "011101110000",
    3145 => "011101101110",
    3146 => "011101101100",
    3147 => "011101101010",
    3148 => "011101101000",
    3149 => "011101100110",
    3150 => "011101100100",
    3151 => "011101100010",
    3152 => "011101100000",
    3153 => "011101011110",
    3154 => "011101011100",
    3155 => "011101011010",
    3156 => "011101011000",
    3157 => "011101010110",
    3158 => "011101010100",
    3159 => "011101010010",
    3160 => "011101010000",
    3161 => "011101001110",
    3162 => "011101001100",
    3163 => "011101001010",
    3164 => "011101001000",
    3165 => "011101000110",
    3166 => "011101000100",
    3167 => "011101000010",
    3168 => "011101000000",
    3169 => "011100111110",
    3170 => "011100111100",
    3171 => "011100111010",
    3172 => "011100111000",
    3173 => "011100110110",
    3174 => "011100110100",
    3175 => "011100110010",
    3176 => "011100110000",
    3177 => "011100101110",
    3178 => "011100101100",
    3179 => "011100101010",
    3180 => "011100101000",
    3181 => "011100100110",
    3182 => "011100100100",
    3183 => "011100100010",
    3184 => "011100100000",
    3185 => "011100011110",
    3186 => "011100011100",
    3187 => "011100011010",
    3188 => "011100011000",
    3189 => "011100010110",
    3190 => "011100010100",
    3191 => "011100010010",
    3192 => "011100010000",
    3193 => "011100001110",
    3194 => "011100001100",
    3195 => "011100001010",
    3196 => "011100001000",
    3197 => "011100000110",
    3198 => "011100000100",
    3199 => "011100000010",
    3200 => "011100000000",
    3201 => "011011111110",
    3202 => "011011111100",
    3203 => "011011111010",
    3204 => "011011111000",
    3205 => "011011110110",
    3206 => "011011110100",
    3207 => "011011110010",
    3208 => "011011110000",
    3209 => "011011101110",
    3210 => "011011101100",
    3211 => "011011101010",
    3212 => "011011101000",
    3213 => "011011100110",
    3214 => "011011100100",
    3215 => "011011100010",
    3216 => "011011100000",
    3217 => "011011011110",
    3218 => "011011011100",
    3219 => "011011011010",
    3220 => "011011011000",
    3221 => "011011010110",
    3222 => "011011010100",
    3223 => "011011010010",
    3224 => "011011010000",
    3225 => "011011001110",
    3226 => "011011001100",
    3227 => "011011001010",
    3228 => "011011001000",
    3229 => "011011000110",
    3230 => "011011000100",
    3231 => "011011000010",
    3232 => "011011000000",
    3233 => "011010111110",
    3234 => "011010111100",
    3235 => "011010111010",
    3236 => "011010111000",
    3237 => "011010110110",
    3238 => "011010110100",
    3239 => "011010110010",
    3240 => "011010110000",
    3241 => "011010101110",
    3242 => "011010101100",
    3243 => "011010101010",
    3244 => "011010101000",
    3245 => "011010100110",
    3246 => "011010100100",
    3247 => "011010100010",
    3248 => "011010100000",
    3249 => "011010011110",
    3250 => "011010011100",
    3251 => "011010011010",
    3252 => "011010011000",
    3253 => "011010010110",
    3254 => "011010010100",
    3255 => "011010010010",
    3256 => "011010010000",
    3257 => "011010001110",
    3258 => "011010001100",
    3259 => "011010001010",
    3260 => "011010001000",
    3261 => "011010000110",
    3262 => "011010000100",
    3263 => "011010000010",
    3264 => "011010000000",
    3265 => "011001111110",
    3266 => "011001111100",
    3267 => "011001111010",
    3268 => "011001111000",
    3269 => "011001110110",
    3270 => "011001110100",
    3271 => "011001110010",
    3272 => "011001110000",
    3273 => "011001101110",
    3274 => "011001101100",
    3275 => "011001101010",
    3276 => "011001101000",
    3277 => "011001100110",
    3278 => "011001100100",
    3279 => "011001100010",
    3280 => "011001100000",
    3281 => "011001011110",
    3282 => "011001011100",
    3283 => "011001011010",
    3284 => "011001011000",
    3285 => "011001010110",
    3286 => "011001010100",
    3287 => "011001010010",
    3288 => "011001010000",
    3289 => "011001001110",
    3290 => "011001001100",
    3291 => "011001001010",
    3292 => "011001001000",
    3293 => "011001000110",
    3294 => "011001000100",
    3295 => "011001000010",
    3296 => "011001000000",
    3297 => "011000111110",
    3298 => "011000111100",
    3299 => "011000111010",
    3300 => "011000111000",
    3301 => "011000110110",
    3302 => "011000110100",
    3303 => "011000110010",
    3304 => "011000110000",
    3305 => "011000101110",
    3306 => "011000101100",
    3307 => "011000101010",
    3308 => "011000101000",
    3309 => "011000100110",
    3310 => "011000100100",
    3311 => "011000100010",
    3312 => "011000100000",
    3313 => "011000011110",
    3314 => "011000011100",
    3315 => "011000011010",
    3316 => "011000011000",
    3317 => "011000010110",
    3318 => "011000010100",
    3319 => "011000010010",
    3320 => "011000010000",
    3321 => "011000001110",
    3322 => "011000001100",
    3323 => "011000001010",
    3324 => "011000001000",
    3325 => "011000000110",
    3326 => "011000000100",
    3327 => "011000000010",
    3328 => "011000000000",
    3329 => "010111111110",
    3330 => "010111111100",
    3331 => "010111111010",
    3332 => "010111111000",
    3333 => "010111110110",
    3334 => "010111110100",
    3335 => "010111110010",
    3336 => "010111110000",
    3337 => "010111101110",
    3338 => "010111101100",
    3339 => "010111101010",
    3340 => "010111101000",
    3341 => "010111100110",
    3342 => "010111100100",
    3343 => "010111100010",
    3344 => "010111100000",
    3345 => "010111011110",
    3346 => "010111011100",
    3347 => "010111011010",
    3348 => "010111011000",
    3349 => "010111010110",
    3350 => "010111010100",
    3351 => "010111010010",
    3352 => "010111010000",
    3353 => "010111001110",
    3354 => "010111001100",
    3355 => "010111001010",
    3356 => "010111001000",
    3357 => "010111000110",
    3358 => "010111000100",
    3359 => "010111000010",
    3360 => "010111000000",
    3361 => "010110111110",
    3362 => "010110111100",
    3363 => "010110111010",
    3364 => "010110111000",
    3365 => "010110110110",
    3366 => "010110110100",
    3367 => "010110110010",
    3368 => "010110110000",
    3369 => "010110101110",
    3370 => "010110101100",
    3371 => "010110101010",
    3372 => "010110101000",
    3373 => "010110100110",
    3374 => "010110100100",
    3375 => "010110100010",
    3376 => "010110100000",
    3377 => "010110011110",
    3378 => "010110011100",
    3379 => "010110011010",
    3380 => "010110011000",
    3381 => "010110010110",
    3382 => "010110010100",
    3383 => "010110010010",
    3384 => "010110010000",
    3385 => "010110001110",
    3386 => "010110001100",
    3387 => "010110001010",
    3388 => "010110001000",
    3389 => "010110000110",
    3390 => "010110000100",
    3391 => "010110000010",
    3392 => "010110000000",
    3393 => "010101111110",
    3394 => "010101111100",
    3395 => "010101111010",
    3396 => "010101111000",
    3397 => "010101110110",
    3398 => "010101110100",
    3399 => "010101110010",
    3400 => "010101110000",
    3401 => "010101101110",
    3402 => "010101101100",
    3403 => "010101101010",
    3404 => "010101101000",
    3405 => "010101100110",
    3406 => "010101100100",
    3407 => "010101100010",
    3408 => "010101100000",
    3409 => "010101011110",
    3410 => "010101011100",
    3411 => "010101011010",
    3412 => "010101011000",
    3413 => "010101010110",
    3414 => "010101010100",
    3415 => "010101010010",
    3416 => "010101010000",
    3417 => "010101001110",
    3418 => "010101001100",
    3419 => "010101001010",
    3420 => "010101001000",
    3421 => "010101000110",
    3422 => "010101000100",
    3423 => "010101000010",
    3424 => "010101000000",
    3425 => "010100111110",
    3426 => "010100111100",
    3427 => "010100111010",
    3428 => "010100111000",
    3429 => "010100110110",
    3430 => "010100110100",
    3431 => "010100110010",
    3432 => "010100110000",
    3433 => "010100101110",
    3434 => "010100101100",
    3435 => "010100101010",
    3436 => "010100101000",
    3437 => "010100100110",
    3438 => "010100100100",
    3439 => "010100100010",
    3440 => "010100100000",
    3441 => "010100011110",
    3442 => "010100011100",
    3443 => "010100011010",
    3444 => "010100011000",
    3445 => "010100010110",
    3446 => "010100010100",
    3447 => "010100010010",
    3448 => "010100010000",
    3449 => "010100001110",
    3450 => "010100001100",
    3451 => "010100001010",
    3452 => "010100001000",
    3453 => "010100000110",
    3454 => "010100000100",
    3455 => "010100000010",
    3456 => "010100000000",
    3457 => "010011111110",
    3458 => "010011111100",
    3459 => "010011111010",
    3460 => "010011111000",
    3461 => "010011110110",
    3462 => "010011110100",
    3463 => "010011110010",
    3464 => "010011110000",
    3465 => "010011101110",
    3466 => "010011101100",
    3467 => "010011101010",
    3468 => "010011101000",
    3469 => "010011100110",
    3470 => "010011100100",
    3471 => "010011100010",
    3472 => "010011100000",
    3473 => "010011011110",
    3474 => "010011011100",
    3475 => "010011011010",
    3476 => "010011011000",
    3477 => "010011010110",
    3478 => "010011010100",
    3479 => "010011010010",
    3480 => "010011010000",
    3481 => "010011001110",
    3482 => "010011001100",
    3483 => "010011001010",
    3484 => "010011001000",
    3485 => "010011000110",
    3486 => "010011000100",
    3487 => "010011000010",
    3488 => "010011000000",
    3489 => "010010111110",
    3490 => "010010111100",
    3491 => "010010111010",
    3492 => "010010111000",
    3493 => "010010110110",
    3494 => "010010110100",
    3495 => "010010110010",
    3496 => "010010110000",
    3497 => "010010101110",
    3498 => "010010101100",
    3499 => "010010101010",
    3500 => "010010101000",
    3501 => "010010100110",
    3502 => "010010100100",
    3503 => "010010100010",
    3504 => "010010100000",
    3505 => "010010011110",
    3506 => "010010011100",
    3507 => "010010011010",
    3508 => "010010011000",
    3509 => "010010010110",
    3510 => "010010010100",
    3511 => "010010010010",
    3512 => "010010010000",
    3513 => "010010001110",
    3514 => "010010001100",
    3515 => "010010001010",
    3516 => "010010001000",
    3517 => "010010000110",
    3518 => "010010000100",
    3519 => "010010000010",
    3520 => "010010000000",
    3521 => "010001111110",
    3522 => "010001111100",
    3523 => "010001111010",
    3524 => "010001111000",
    3525 => "010001110110",
    3526 => "010001110100",
    3527 => "010001110010",
    3528 => "010001110000",
    3529 => "010001101110",
    3530 => "010001101100",
    3531 => "010001101010",
    3532 => "010001101000",
    3533 => "010001100110",
    3534 => "010001100100",
    3535 => "010001100010",
    3536 => "010001100000",
    3537 => "010001011110",
    3538 => "010001011100",
    3539 => "010001011010",
    3540 => "010001011000",
    3541 => "010001010110",
    3542 => "010001010100",
    3543 => "010001010010",
    3544 => "010001010000",
    3545 => "010001001110",
    3546 => "010001001100",
    3547 => "010001001010",
    3548 => "010001001000",
    3549 => "010001000110",
    3550 => "010001000100",
    3551 => "010001000010",
    3552 => "010001000000",
    3553 => "010000111110",
    3554 => "010000111100",
    3555 => "010000111010",
    3556 => "010000111000",
    3557 => "010000110110",
    3558 => "010000110100",
    3559 => "010000110010",
    3560 => "010000110000",
    3561 => "010000101110",
    3562 => "010000101100",
    3563 => "010000101010",
    3564 => "010000101000",
    3565 => "010000100110",
    3566 => "010000100100",
    3567 => "010000100010",
    3568 => "010000100000",
    3569 => "010000011110",
    3570 => "010000011100",
    3571 => "010000011010",
    3572 => "010000011000",
    3573 => "010000010110",
    3574 => "010000010100",
    3575 => "010000010010",
    3576 => "010000010000",
    3577 => "010000001110",
    3578 => "010000001100",
    3579 => "010000001010",
    3580 => "010000001000",
    3581 => "010000000110",
    3582 => "010000000100",
    3583 => "010000000010",
    3584 => "010000000000",
    3585 => "001111111110",
    3586 => "001111111100",
    3587 => "001111111010",
    3588 => "001111111000",
    3589 => "001111110110",
    3590 => "001111110100",
    3591 => "001111110010",
    3592 => "001111110000",
    3593 => "001111101110",
    3594 => "001111101100",
    3595 => "001111101010",
    3596 => "001111101000",
    3597 => "001111100110",
    3598 => "001111100100",
    3599 => "001111100010",
    3600 => "001111100000",
    3601 => "001111011110",
    3602 => "001111011100",
    3603 => "001111011010",
    3604 => "001111011000",
    3605 => "001111010110",
    3606 => "001111010100",
    3607 => "001111010010",
    3608 => "001111010000",
    3609 => "001111001110",
    3610 => "001111001100",
    3611 => "001111001010",
    3612 => "001111001000",
    3613 => "001111000110",
    3614 => "001111000100",
    3615 => "001111000010",
    3616 => "001111000000",
    3617 => "001110111110",
    3618 => "001110111100",
    3619 => "001110111010",
    3620 => "001110111000",
    3621 => "001110110110",
    3622 => "001110110100",
    3623 => "001110110010",
    3624 => "001110110000",
    3625 => "001110101110",
    3626 => "001110101100",
    3627 => "001110101010",
    3628 => "001110101000",
    3629 => "001110100110",
    3630 => "001110100100",
    3631 => "001110100010",
    3632 => "001110100000",
    3633 => "001110011110",
    3634 => "001110011100",
    3635 => "001110011010",
    3636 => "001110011000",
    3637 => "001110010110",
    3638 => "001110010100",
    3639 => "001110010010",
    3640 => "001110010000",
    3641 => "001110001110",
    3642 => "001110001100",
    3643 => "001110001010",
    3644 => "001110001000",
    3645 => "001110000110",
    3646 => "001110000100",
    3647 => "001110000010",
    3648 => "001110000000",
    3649 => "001101111110",
    3650 => "001101111100",
    3651 => "001101111010",
    3652 => "001101111000",
    3653 => "001101110110",
    3654 => "001101110100",
    3655 => "001101110010",
    3656 => "001101110000",
    3657 => "001101101110",
    3658 => "001101101100",
    3659 => "001101101010",
    3660 => "001101101000",
    3661 => "001101100110",
    3662 => "001101100100",
    3663 => "001101100010",
    3664 => "001101100000",
    3665 => "001101011110",
    3666 => "001101011100",
    3667 => "001101011010",
    3668 => "001101011000",
    3669 => "001101010110",
    3670 => "001101010100",
    3671 => "001101010010",
    3672 => "001101010000",
    3673 => "001101001110",
    3674 => "001101001100",
    3675 => "001101001010",
    3676 => "001101001000",
    3677 => "001101000110",
    3678 => "001101000100",
    3679 => "001101000010",
    3680 => "001101000000",
    3681 => "001100111110",
    3682 => "001100111100",
    3683 => "001100111010",
    3684 => "001100111000",
    3685 => "001100110110",
    3686 => "001100110100",
    3687 => "001100110010",
    3688 => "001100110000",
    3689 => "001100101110",
    3690 => "001100101100",
    3691 => "001100101010",
    3692 => "001100101000",
    3693 => "001100100110",
    3694 => "001100100100",
    3695 => "001100100010",
    3696 => "001100100000",
    3697 => "001100011110",
    3698 => "001100011100",
    3699 => "001100011010",
    3700 => "001100011000",
    3701 => "001100010110",
    3702 => "001100010100",
    3703 => "001100010010",
    3704 => "001100010000",
    3705 => "001100001110",
    3706 => "001100001100",
    3707 => "001100001010",
    3708 => "001100001000",
    3709 => "001100000110",
    3710 => "001100000100",
    3711 => "001100000010",
    3712 => "001100000000",
    3713 => "001011111110",
    3714 => "001011111100",
    3715 => "001011111010",
    3716 => "001011111000",
    3717 => "001011110110",
    3718 => "001011110100",
    3719 => "001011110010",
    3720 => "001011110000",
    3721 => "001011101110",
    3722 => "001011101100",
    3723 => "001011101010",
    3724 => "001011101000",
    3725 => "001011100110",
    3726 => "001011100100",
    3727 => "001011100010",
    3728 => "001011100000",
    3729 => "001011011110",
    3730 => "001011011100",
    3731 => "001011011010",
    3732 => "001011011000",
    3733 => "001011010110",
    3734 => "001011010100",
    3735 => "001011010010",
    3736 => "001011010000",
    3737 => "001011001110",
    3738 => "001011001100",
    3739 => "001011001010",
    3740 => "001011001000",
    3741 => "001011000110",
    3742 => "001011000100",
    3743 => "001011000010",
    3744 => "001011000000",
    3745 => "001010111110",
    3746 => "001010111100",
    3747 => "001010111010",
    3748 => "001010111000",
    3749 => "001010110110",
    3750 => "001010110100",
    3751 => "001010110010",
    3752 => "001010110000",
    3753 => "001010101110",
    3754 => "001010101100",
    3755 => "001010101010",
    3756 => "001010101000",
    3757 => "001010100110",
    3758 => "001010100100",
    3759 => "001010100010",
    3760 => "001010100000",
    3761 => "001010011110",
    3762 => "001010011100",
    3763 => "001010011010",
    3764 => "001010011000",
    3765 => "001010010110",
    3766 => "001010010100",
    3767 => "001010010010",
    3768 => "001010010000",
    3769 => "001010001110",
    3770 => "001010001100",
    3771 => "001010001010",
    3772 => "001010001000",
    3773 => "001010000110",
    3774 => "001010000100",
    3775 => "001010000010",
    3776 => "001010000000",
    3777 => "001001111110",
    3778 => "001001111100",
    3779 => "001001111010",
    3780 => "001001111000",
    3781 => "001001110110",
    3782 => "001001110100",
    3783 => "001001110010",
    3784 => "001001110000",
    3785 => "001001101110",
    3786 => "001001101100",
    3787 => "001001101010",
    3788 => "001001101000",
    3789 => "001001100110",
    3790 => "001001100100",
    3791 => "001001100010",
    3792 => "001001100000",
    3793 => "001001011110",
    3794 => "001001011100",
    3795 => "001001011010",
    3796 => "001001011000",
    3797 => "001001010110",
    3798 => "001001010100",
    3799 => "001001010010",
    3800 => "001001010000",
    3801 => "001001001110",
    3802 => "001001001100",
    3803 => "001001001010",
    3804 => "001001001000",
    3805 => "001001000110",
    3806 => "001001000100",
    3807 => "001001000010",
    3808 => "001001000000",
    3809 => "001000111110",
    3810 => "001000111100",
    3811 => "001000111010",
    3812 => "001000111000",
    3813 => "001000110110",
    3814 => "001000110100",
    3815 => "001000110010",
    3816 => "001000110000",
    3817 => "001000101110",
    3818 => "001000101100",
    3819 => "001000101010",
    3820 => "001000101000",
    3821 => "001000100110",
    3822 => "001000100100",
    3823 => "001000100010",
    3824 => "001000100000",
    3825 => "001000011110",
    3826 => "001000011100",
    3827 => "001000011010",
    3828 => "001000011000",
    3829 => "001000010110",
    3830 => "001000010100",
    3831 => "001000010010",
    3832 => "001000010000",
    3833 => "001000001110",
    3834 => "001000001100",
    3835 => "001000001010",
    3836 => "001000001000",
    3837 => "001000000110",
    3838 => "001000000100",
    3839 => "001000000010",
    3840 => "001000000000",
    3841 => "000111111110",
    3842 => "000111111100",
    3843 => "000111111010",
    3844 => "000111111000",
    3845 => "000111110110",
    3846 => "000111110100",
    3847 => "000111110010",
    3848 => "000111110000",
    3849 => "000111101110",
    3850 => "000111101100",
    3851 => "000111101010",
    3852 => "000111101000",
    3853 => "000111100110",
    3854 => "000111100100",
    3855 => "000111100010",
    3856 => "000111100000",
    3857 => "000111011110",
    3858 => "000111011100",
    3859 => "000111011010",
    3860 => "000111011000",
    3861 => "000111010110",
    3862 => "000111010100",
    3863 => "000111010010",
    3864 => "000111010000",
    3865 => "000111001110",
    3866 => "000111001100",
    3867 => "000111001010",
    3868 => "000111001000",
    3869 => "000111000110",
    3870 => "000111000100",
    3871 => "000111000010",
    3872 => "000111000000",
    3873 => "000110111110",
    3874 => "000110111100",
    3875 => "000110111010",
    3876 => "000110111000",
    3877 => "000110110110",
    3878 => "000110110100",
    3879 => "000110110010",
    3880 => "000110110000",
    3881 => "000110101110",
    3882 => "000110101100",
    3883 => "000110101010",
    3884 => "000110101000",
    3885 => "000110100110",
    3886 => "000110100100",
    3887 => "000110100010",
    3888 => "000110100000",
    3889 => "000110011110",
    3890 => "000110011100",
    3891 => "000110011010",
    3892 => "000110011000",
    3893 => "000110010110",
    3894 => "000110010100",
    3895 => "000110010010",
    3896 => "000110010000",
    3897 => "000110001110",
    3898 => "000110001100",
    3899 => "000110001010",
    3900 => "000110001000",
    3901 => "000110000110",
    3902 => "000110000100",
    3903 => "000110000010",
    3904 => "000110000000",
    3905 => "000101111110",
    3906 => "000101111100",
    3907 => "000101111010",
    3908 => "000101111000",
    3909 => "000101110110",
    3910 => "000101110100",
    3911 => "000101110010",
    3912 => "000101110000",
    3913 => "000101101110",
    3914 => "000101101100",
    3915 => "000101101010",
    3916 => "000101101000",
    3917 => "000101100110",
    3918 => "000101100100",
    3919 => "000101100010",
    3920 => "000101100000",
    3921 => "000101011110",
    3922 => "000101011100",
    3923 => "000101011010",
    3924 => "000101011000",
    3925 => "000101010110",
    3926 => "000101010100",
    3927 => "000101010010",
    3928 => "000101010000",
    3929 => "000101001110",
    3930 => "000101001100",
    3931 => "000101001010",
    3932 => "000101001000",
    3933 => "000101000110",
    3934 => "000101000100",
    3935 => "000101000010",
    3936 => "000101000000",
    3937 => "000100111110",
    3938 => "000100111100",
    3939 => "000100111010",
    3940 => "000100111000",
    3941 => "000100110110",
    3942 => "000100110100",
    3943 => "000100110010",
    3944 => "000100110000",
    3945 => "000100101110",
    3946 => "000100101100",
    3947 => "000100101010",
    3948 => "000100101000",
    3949 => "000100100110",
    3950 => "000100100100",
    3951 => "000100100010",
    3952 => "000100100000",
    3953 => "000100011110",
    3954 => "000100011100",
    3955 => "000100011010",
    3956 => "000100011000",
    3957 => "000100010110",
    3958 => "000100010100",
    3959 => "000100010010",
    3960 => "000100010000",
    3961 => "000100001110",
    3962 => "000100001100",
    3963 => "000100001010",
    3964 => "000100001000",
    3965 => "000100000110",
    3966 => "000100000100",
    3967 => "000100000010",
    3968 => "000100000000",
    3969 => "000011111110",
    3970 => "000011111100",
    3971 => "000011111010",
    3972 => "000011111000",
    3973 => "000011110110",
    3974 => "000011110100",
    3975 => "000011110010",
    3976 => "000011110000",
    3977 => "000011101110",
    3978 => "000011101100",
    3979 => "000011101010",
    3980 => "000011101000",
    3981 => "000011100110",
    3982 => "000011100100",
    3983 => "000011100010",
    3984 => "000011100000",
    3985 => "000011011110",
    3986 => "000011011100",
    3987 => "000011011010",
    3988 => "000011011000",
    3989 => "000011010110",
    3990 => "000011010100",
    3991 => "000011010010",
    3992 => "000011010000",
    3993 => "000011001110",
    3994 => "000011001100",
    3995 => "000011001010",
    3996 => "000011001000",
    3997 => "000011000110",
    3998 => "000011000100",
    3999 => "000011000010",
    4000 => "000011000000",
    4001 => "000010111110",
    4002 => "000010111100",
    4003 => "000010111010",
    4004 => "000010111000",
    4005 => "000010110110",
    4006 => "000010110100",
    4007 => "000010110010",
    4008 => "000010110000",
    4009 => "000010101110",
    4010 => "000010101100",
    4011 => "000010101010",
    4012 => "000010101000",
    4013 => "000010100110",
    4014 => "000010100100",
    4015 => "000010100010",
    4016 => "000010100000",
    4017 => "000010011110",
    4018 => "000010011100",
    4019 => "000010011010",
    4020 => "000010011000",
    4021 => "000010010110",
    4022 => "000010010100",
    4023 => "000010010010",
    4024 => "000010010000",
    4025 => "000010001110",
    4026 => "000010001100",
    4027 => "000010001010",
    4028 => "000010001000",
    4029 => "000010000110",
    4030 => "000010000100",
    4031 => "000010000010",
    4032 => "000010000000",
    4033 => "000001111110",
    4034 => "000001111100",
    4035 => "000001111010",
    4036 => "000001111000",
    4037 => "000001110110",
    4038 => "000001110100",
    4039 => "000001110010",
    4040 => "000001110000",
    4041 => "000001101110",
    4042 => "000001101100",
    4043 => "000001101010",
    4044 => "000001101000",
    4045 => "000001100110",
    4046 => "000001100100",
    4047 => "000001100010",
    4048 => "000001100000",
    4049 => "000001011110",
    4050 => "000001011100",
    4051 => "000001011010",
    4052 => "000001011000",
    4053 => "000001010110",
    4054 => "000001010100",
    4055 => "000001010010",
    4056 => "000001010000",
    4057 => "000001001110",
    4058 => "000001001100",
    4059 => "000001001010",
    4060 => "000001001000",
    4061 => "000001000110",
    4062 => "000001000100",
    4063 => "000001000010",
    4064 => "000001000000",
    4065 => "000000111110",
    4066 => "000000111100",
    4067 => "000000111010",
    4068 => "000000111000",
    4069 => "000000110110",
    4070 => "000000110100",
    4071 => "000000110010",
    4072 => "000000110000",
    4073 => "000000101110",
    4074 => "000000101100",
    4075 => "000000101010",
    4076 => "000000101000",
    4077 => "000000100110",
    4078 => "000000100100",
    4079 => "000000100010",
    4080 => "000000100000",
    4081 => "000000011110",
    4082 => "000000011100",
    4083 => "000000011010",
    4084 => "000000011000",
    4085 => "000000010110",
    4086 => "000000010100",
    4087 => "000000010010",
    4088 => "000000010000",
    4089 => "000000001110",
    4090 => "000000001100",
    4091 => "000000001010",
    4092 => "000000001000",
    4093 => "000000000110",
    4094 => "000000000100",
    4095 => "000000000100");
begin
 process (address)
 begin
  case address is
     when "000000000000" => data <= triangle_rom(0);
     when "000000000001" => data <= triangle_rom(1);
     when "000000000010" => data <= triangle_rom(2);
     when "000000000011" => data <= triangle_rom(3);
     when "000000000100" => data <= triangle_rom(4);
     when "000000000101" => data <= triangle_rom(5);
     when "000000000110" => data <= triangle_rom(6);
     when "000000000111" => data <= triangle_rom(7);
     when "000000001000" => data <= triangle_rom(8);
     when "000000001001" => data <= triangle_rom(9);
     when "000000001010" => data <= triangle_rom(10);
     when "000000001011" => data <= triangle_rom(11);
     when "000000001100" => data <= triangle_rom(12);
     when "000000001101" => data <= triangle_rom(13);
     when "000000001110" => data <= triangle_rom(14);
     when "000000001111" => data <= triangle_rom(15);
     when "000000010000" => data <= triangle_rom(16);
     when "000000010001" => data <= triangle_rom(17);
     when "000000010010" => data <= triangle_rom(18);
     when "000000010011" => data <= triangle_rom(19);
     when "000000010100" => data <= triangle_rom(20);
     when "000000010101" => data <= triangle_rom(21);
     when "000000010110" => data <= triangle_rom(22);
     when "000000010111" => data <= triangle_rom(23);
     when "000000011000" => data <= triangle_rom(24);
     when "000000011001" => data <= triangle_rom(25);
     when "000000011010" => data <= triangle_rom(26);
     when "000000011011" => data <= triangle_rom(27);
     when "000000011100" => data <= triangle_rom(28);
     when "000000011101" => data <= triangle_rom(29);
     when "000000011110" => data <= triangle_rom(30);
     when "000000011111" => data <= triangle_rom(31);
     when "000000100000" => data <= triangle_rom(32);
     when "000000100001" => data <= triangle_rom(33);
     when "000000100010" => data <= triangle_rom(34);
     when "000000100011" => data <= triangle_rom(35);
     when "000000100100" => data <= triangle_rom(36);
     when "000000100101" => data <= triangle_rom(37);
     when "000000100110" => data <= triangle_rom(38);
     when "000000100111" => data <= triangle_rom(39);
     when "000000101000" => data <= triangle_rom(40);
     when "000000101001" => data <= triangle_rom(41);
     when "000000101010" => data <= triangle_rom(42);
     when "000000101011" => data <= triangle_rom(43);
     when "000000101100" => data <= triangle_rom(44);
     when "000000101101" => data <= triangle_rom(45);
     when "000000101110" => data <= triangle_rom(46);
     when "000000101111" => data <= triangle_rom(47);
     when "000000110000" => data <= triangle_rom(48);
     when "000000110001" => data <= triangle_rom(49);
     when "000000110010" => data <= triangle_rom(50);
     when "000000110011" => data <= triangle_rom(51);
     when "000000110100" => data <= triangle_rom(52);
     when "000000110101" => data <= triangle_rom(53);
     when "000000110110" => data <= triangle_rom(54);
     when "000000110111" => data <= triangle_rom(55);
     when "000000111000" => data <= triangle_rom(56);
     when "000000111001" => data <= triangle_rom(57);
     when "000000111010" => data <= triangle_rom(58);
     when "000000111011" => data <= triangle_rom(59);
     when "000000111100" => data <= triangle_rom(60);
     when "000000111101" => data <= triangle_rom(61);
     when "000000111110" => data <= triangle_rom(62);
     when "000000111111" => data <= triangle_rom(63);
     when "000001000000" => data <= triangle_rom(64);
     when "000001000001" => data <= triangle_rom(65);
     when "000001000010" => data <= triangle_rom(66);
     when "000001000011" => data <= triangle_rom(67);
     when "000001000100" => data <= triangle_rom(68);
     when "000001000101" => data <= triangle_rom(69);
     when "000001000110" => data <= triangle_rom(70);
     when "000001000111" => data <= triangle_rom(71);
     when "000001001000" => data <= triangle_rom(72);
     when "000001001001" => data <= triangle_rom(73);
     when "000001001010" => data <= triangle_rom(74);
     when "000001001011" => data <= triangle_rom(75);
     when "000001001100" => data <= triangle_rom(76);
     when "000001001101" => data <= triangle_rom(77);
     when "000001001110" => data <= triangle_rom(78);
     when "000001001111" => data <= triangle_rom(79);
     when "000001010000" => data <= triangle_rom(80);
     when "000001010001" => data <= triangle_rom(81);
     when "000001010010" => data <= triangle_rom(82);
     when "000001010011" => data <= triangle_rom(83);
     when "000001010100" => data <= triangle_rom(84);
     when "000001010101" => data <= triangle_rom(85);
     when "000001010110" => data <= triangle_rom(86);
     when "000001010111" => data <= triangle_rom(87);
     when "000001011000" => data <= triangle_rom(88);
     when "000001011001" => data <= triangle_rom(89);
     when "000001011010" => data <= triangle_rom(90);
     when "000001011011" => data <= triangle_rom(91);
     when "000001011100" => data <= triangle_rom(92);
     when "000001011101" => data <= triangle_rom(93);
     when "000001011110" => data <= triangle_rom(94);
     when "000001011111" => data <= triangle_rom(95);
     when "000001100000" => data <= triangle_rom(96);
     when "000001100001" => data <= triangle_rom(97);
     when "000001100010" => data <= triangle_rom(98);
     when "000001100011" => data <= triangle_rom(99);
     when "000001100100" => data <= triangle_rom(100);
     when "000001100101" => data <= triangle_rom(101);
     when "000001100110" => data <= triangle_rom(102);
     when "000001100111" => data <= triangle_rom(103);
     when "000001101000" => data <= triangle_rom(104);
     when "000001101001" => data <= triangle_rom(105);
     when "000001101010" => data <= triangle_rom(106);
     when "000001101011" => data <= triangle_rom(107);
     when "000001101100" => data <= triangle_rom(108);
     when "000001101101" => data <= triangle_rom(109);
     when "000001101110" => data <= triangle_rom(110);
     when "000001101111" => data <= triangle_rom(111);
     when "000001110000" => data <= triangle_rom(112);
     when "000001110001" => data <= triangle_rom(113);
     when "000001110010" => data <= triangle_rom(114);
     when "000001110011" => data <= triangle_rom(115);
     when "000001110100" => data <= triangle_rom(116);
     when "000001110101" => data <= triangle_rom(117);
     when "000001110110" => data <= triangle_rom(118);
     when "000001110111" => data <= triangle_rom(119);
     when "000001111000" => data <= triangle_rom(120);
     when "000001111001" => data <= triangle_rom(121);
     when "000001111010" => data <= triangle_rom(122);
     when "000001111011" => data <= triangle_rom(123);
     when "000001111100" => data <= triangle_rom(124);
     when "000001111101" => data <= triangle_rom(125);
     when "000001111110" => data <= triangle_rom(126);
     when "000001111111" => data <= triangle_rom(127);
     when "000010000000" => data <= triangle_rom(128);
     when "000010000001" => data <= triangle_rom(129);
     when "000010000010" => data <= triangle_rom(130);
     when "000010000011" => data <= triangle_rom(131);
     when "000010000100" => data <= triangle_rom(132);
     when "000010000101" => data <= triangle_rom(133);
     when "000010000110" => data <= triangle_rom(134);
     when "000010000111" => data <= triangle_rom(135);
     when "000010001000" => data <= triangle_rom(136);
     when "000010001001" => data <= triangle_rom(137);
     when "000010001010" => data <= triangle_rom(138);
     when "000010001011" => data <= triangle_rom(139);
     when "000010001100" => data <= triangle_rom(140);
     when "000010001101" => data <= triangle_rom(141);
     when "000010001110" => data <= triangle_rom(142);
     when "000010001111" => data <= triangle_rom(143);
     when "000010010000" => data <= triangle_rom(144);
     when "000010010001" => data <= triangle_rom(145);
     when "000010010010" => data <= triangle_rom(146);
     when "000010010011" => data <= triangle_rom(147);
     when "000010010100" => data <= triangle_rom(148);
     when "000010010101" => data <= triangle_rom(149);
     when "000010010110" => data <= triangle_rom(150);
     when "000010010111" => data <= triangle_rom(151);
     when "000010011000" => data <= triangle_rom(152);
     when "000010011001" => data <= triangle_rom(153);
     when "000010011010" => data <= triangle_rom(154);
     when "000010011011" => data <= triangle_rom(155);
     when "000010011100" => data <= triangle_rom(156);
     when "000010011101" => data <= triangle_rom(157);
     when "000010011110" => data <= triangle_rom(158);
     when "000010011111" => data <= triangle_rom(159);
     when "000010100000" => data <= triangle_rom(160);
     when "000010100001" => data <= triangle_rom(161);
     when "000010100010" => data <= triangle_rom(162);
     when "000010100011" => data <= triangle_rom(163);
     when "000010100100" => data <= triangle_rom(164);
     when "000010100101" => data <= triangle_rom(165);
     when "000010100110" => data <= triangle_rom(166);
     when "000010100111" => data <= triangle_rom(167);
     when "000010101000" => data <= triangle_rom(168);
     when "000010101001" => data <= triangle_rom(169);
     when "000010101010" => data <= triangle_rom(170);
     when "000010101011" => data <= triangle_rom(171);
     when "000010101100" => data <= triangle_rom(172);
     when "000010101101" => data <= triangle_rom(173);
     when "000010101110" => data <= triangle_rom(174);
     when "000010101111" => data <= triangle_rom(175);
     when "000010110000" => data <= triangle_rom(176);
     when "000010110001" => data <= triangle_rom(177);
     when "000010110010" => data <= triangle_rom(178);
     when "000010110011" => data <= triangle_rom(179);
     when "000010110100" => data <= triangle_rom(180);
     when "000010110101" => data <= triangle_rom(181);
     when "000010110110" => data <= triangle_rom(182);
     when "000010110111" => data <= triangle_rom(183);
     when "000010111000" => data <= triangle_rom(184);
     when "000010111001" => data <= triangle_rom(185);
     when "000010111010" => data <= triangle_rom(186);
     when "000010111011" => data <= triangle_rom(187);
     when "000010111100" => data <= triangle_rom(188);
     when "000010111101" => data <= triangle_rom(189);
     when "000010111110" => data <= triangle_rom(190);
     when "000010111111" => data <= triangle_rom(191);
     when "000011000000" => data <= triangle_rom(192);
     when "000011000001" => data <= triangle_rom(193);
     when "000011000010" => data <= triangle_rom(194);
     when "000011000011" => data <= triangle_rom(195);
     when "000011000100" => data <= triangle_rom(196);
     when "000011000101" => data <= triangle_rom(197);
     when "000011000110" => data <= triangle_rom(198);
     when "000011000111" => data <= triangle_rom(199);
     when "000011001000" => data <= triangle_rom(200);
     when "000011001001" => data <= triangle_rom(201);
     when "000011001010" => data <= triangle_rom(202);
     when "000011001011" => data <= triangle_rom(203);
     when "000011001100" => data <= triangle_rom(204);
     when "000011001101" => data <= triangle_rom(205);
     when "000011001110" => data <= triangle_rom(206);
     when "000011001111" => data <= triangle_rom(207);
     when "000011010000" => data <= triangle_rom(208);
     when "000011010001" => data <= triangle_rom(209);
     when "000011010010" => data <= triangle_rom(210);
     when "000011010011" => data <= triangle_rom(211);
     when "000011010100" => data <= triangle_rom(212);
     when "000011010101" => data <= triangle_rom(213);
     when "000011010110" => data <= triangle_rom(214);
     when "000011010111" => data <= triangle_rom(215);
     when "000011011000" => data <= triangle_rom(216);
     when "000011011001" => data <= triangle_rom(217);
     when "000011011010" => data <= triangle_rom(218);
     when "000011011011" => data <= triangle_rom(219);
     when "000011011100" => data <= triangle_rom(220);
     when "000011011101" => data <= triangle_rom(221);
     when "000011011110" => data <= triangle_rom(222);
     when "000011011111" => data <= triangle_rom(223);
     when "000011100000" => data <= triangle_rom(224);
     when "000011100001" => data <= triangle_rom(225);
     when "000011100010" => data <= triangle_rom(226);
     when "000011100011" => data <= triangle_rom(227);
     when "000011100100" => data <= triangle_rom(228);
     when "000011100101" => data <= triangle_rom(229);
     when "000011100110" => data <= triangle_rom(230);
     when "000011100111" => data <= triangle_rom(231);
     when "000011101000" => data <= triangle_rom(232);
     when "000011101001" => data <= triangle_rom(233);
     when "000011101010" => data <= triangle_rom(234);
     when "000011101011" => data <= triangle_rom(235);
     when "000011101100" => data <= triangle_rom(236);
     when "000011101101" => data <= triangle_rom(237);
     when "000011101110" => data <= triangle_rom(238);
     when "000011101111" => data <= triangle_rom(239);
     when "000011110000" => data <= triangle_rom(240);
     when "000011110001" => data <= triangle_rom(241);
     when "000011110010" => data <= triangle_rom(242);
     when "000011110011" => data <= triangle_rom(243);
     when "000011110100" => data <= triangle_rom(244);
     when "000011110101" => data <= triangle_rom(245);
     when "000011110110" => data <= triangle_rom(246);
     when "000011110111" => data <= triangle_rom(247);
     when "000011111000" => data <= triangle_rom(248);
     when "000011111001" => data <= triangle_rom(249);
     when "000011111010" => data <= triangle_rom(250);
     when "000011111011" => data <= triangle_rom(251);
     when "000011111100" => data <= triangle_rom(252);
     when "000011111101" => data <= triangle_rom(253);
     when "000011111110" => data <= triangle_rom(254);
     when "000011111111" => data <= triangle_rom(255);
     when "000100000000" => data <= triangle_rom(256);
     when "000100000001" => data <= triangle_rom(257);
     when "000100000010" => data <= triangle_rom(258);
     when "000100000011" => data <= triangle_rom(259);
     when "000100000100" => data <= triangle_rom(260);
     when "000100000101" => data <= triangle_rom(261);
     when "000100000110" => data <= triangle_rom(262);
     when "000100000111" => data <= triangle_rom(263);
     when "000100001000" => data <= triangle_rom(264);
     when "000100001001" => data <= triangle_rom(265);
     when "000100001010" => data <= triangle_rom(266);
     when "000100001011" => data <= triangle_rom(267);
     when "000100001100" => data <= triangle_rom(268);
     when "000100001101" => data <= triangle_rom(269);
     when "000100001110" => data <= triangle_rom(270);
     when "000100001111" => data <= triangle_rom(271);
     when "000100010000" => data <= triangle_rom(272);
     when "000100010001" => data <= triangle_rom(273);
     when "000100010010" => data <= triangle_rom(274);
     when "000100010011" => data <= triangle_rom(275);
     when "000100010100" => data <= triangle_rom(276);
     when "000100010101" => data <= triangle_rom(277);
     when "000100010110" => data <= triangle_rom(278);
     when "000100010111" => data <= triangle_rom(279);
     when "000100011000" => data <= triangle_rom(280);
     when "000100011001" => data <= triangle_rom(281);
     when "000100011010" => data <= triangle_rom(282);
     when "000100011011" => data <= triangle_rom(283);
     when "000100011100" => data <= triangle_rom(284);
     when "000100011101" => data <= triangle_rom(285);
     when "000100011110" => data <= triangle_rom(286);
     when "000100011111" => data <= triangle_rom(287);
     when "000100100000" => data <= triangle_rom(288);
     when "000100100001" => data <= triangle_rom(289);
     when "000100100010" => data <= triangle_rom(290);
     when "000100100011" => data <= triangle_rom(291);
     when "000100100100" => data <= triangle_rom(292);
     when "000100100101" => data <= triangle_rom(293);
     when "000100100110" => data <= triangle_rom(294);
     when "000100100111" => data <= triangle_rom(295);
     when "000100101000" => data <= triangle_rom(296);
     when "000100101001" => data <= triangle_rom(297);
     when "000100101010" => data <= triangle_rom(298);
     when "000100101011" => data <= triangle_rom(299);
     when "000100101100" => data <= triangle_rom(300);
     when "000100101101" => data <= triangle_rom(301);
     when "000100101110" => data <= triangle_rom(302);
     when "000100101111" => data <= triangle_rom(303);
     when "000100110000" => data <= triangle_rom(304);
     when "000100110001" => data <= triangle_rom(305);
     when "000100110010" => data <= triangle_rom(306);
     when "000100110011" => data <= triangle_rom(307);
     when "000100110100" => data <= triangle_rom(308);
     when "000100110101" => data <= triangle_rom(309);
     when "000100110110" => data <= triangle_rom(310);
     when "000100110111" => data <= triangle_rom(311);
     when "000100111000" => data <= triangle_rom(312);
     when "000100111001" => data <= triangle_rom(313);
     when "000100111010" => data <= triangle_rom(314);
     when "000100111011" => data <= triangle_rom(315);
     when "000100111100" => data <= triangle_rom(316);
     when "000100111101" => data <= triangle_rom(317);
     when "000100111110" => data <= triangle_rom(318);
     when "000100111111" => data <= triangle_rom(319);
     when "000101000000" => data <= triangle_rom(320);
     when "000101000001" => data <= triangle_rom(321);
     when "000101000010" => data <= triangle_rom(322);
     when "000101000011" => data <= triangle_rom(323);
     when "000101000100" => data <= triangle_rom(324);
     when "000101000101" => data <= triangle_rom(325);
     when "000101000110" => data <= triangle_rom(326);
     when "000101000111" => data <= triangle_rom(327);
     when "000101001000" => data <= triangle_rom(328);
     when "000101001001" => data <= triangle_rom(329);
     when "000101001010" => data <= triangle_rom(330);
     when "000101001011" => data <= triangle_rom(331);
     when "000101001100" => data <= triangle_rom(332);
     when "000101001101" => data <= triangle_rom(333);
     when "000101001110" => data <= triangle_rom(334);
     when "000101001111" => data <= triangle_rom(335);
     when "000101010000" => data <= triangle_rom(336);
     when "000101010001" => data <= triangle_rom(337);
     when "000101010010" => data <= triangle_rom(338);
     when "000101010011" => data <= triangle_rom(339);
     when "000101010100" => data <= triangle_rom(340);
     when "000101010101" => data <= triangle_rom(341);
     when "000101010110" => data <= triangle_rom(342);
     when "000101010111" => data <= triangle_rom(343);
     when "000101011000" => data <= triangle_rom(344);
     when "000101011001" => data <= triangle_rom(345);
     when "000101011010" => data <= triangle_rom(346);
     when "000101011011" => data <= triangle_rom(347);
     when "000101011100" => data <= triangle_rom(348);
     when "000101011101" => data <= triangle_rom(349);
     when "000101011110" => data <= triangle_rom(350);
     when "000101011111" => data <= triangle_rom(351);
     when "000101100000" => data <= triangle_rom(352);
     when "000101100001" => data <= triangle_rom(353);
     when "000101100010" => data <= triangle_rom(354);
     when "000101100011" => data <= triangle_rom(355);
     when "000101100100" => data <= triangle_rom(356);
     when "000101100101" => data <= triangle_rom(357);
     when "000101100110" => data <= triangle_rom(358);
     when "000101100111" => data <= triangle_rom(359);
     when "000101101000" => data <= triangle_rom(360);
     when "000101101001" => data <= triangle_rom(361);
     when "000101101010" => data <= triangle_rom(362);
     when "000101101011" => data <= triangle_rom(363);
     when "000101101100" => data <= triangle_rom(364);
     when "000101101101" => data <= triangle_rom(365);
     when "000101101110" => data <= triangle_rom(366);
     when "000101101111" => data <= triangle_rom(367);
     when "000101110000" => data <= triangle_rom(368);
     when "000101110001" => data <= triangle_rom(369);
     when "000101110010" => data <= triangle_rom(370);
     when "000101110011" => data <= triangle_rom(371);
     when "000101110100" => data <= triangle_rom(372);
     when "000101110101" => data <= triangle_rom(373);
     when "000101110110" => data <= triangle_rom(374);
     when "000101110111" => data <= triangle_rom(375);
     when "000101111000" => data <= triangle_rom(376);
     when "000101111001" => data <= triangle_rom(377);
     when "000101111010" => data <= triangle_rom(378);
     when "000101111011" => data <= triangle_rom(379);
     when "000101111100" => data <= triangle_rom(380);
     when "000101111101" => data <= triangle_rom(381);
     when "000101111110" => data <= triangle_rom(382);
     when "000101111111" => data <= triangle_rom(383);
     when "000110000000" => data <= triangle_rom(384);
     when "000110000001" => data <= triangle_rom(385);
     when "000110000010" => data <= triangle_rom(386);
     when "000110000011" => data <= triangle_rom(387);
     when "000110000100" => data <= triangle_rom(388);
     when "000110000101" => data <= triangle_rom(389);
     when "000110000110" => data <= triangle_rom(390);
     when "000110000111" => data <= triangle_rom(391);
     when "000110001000" => data <= triangle_rom(392);
     when "000110001001" => data <= triangle_rom(393);
     when "000110001010" => data <= triangle_rom(394);
     when "000110001011" => data <= triangle_rom(395);
     when "000110001100" => data <= triangle_rom(396);
     when "000110001101" => data <= triangle_rom(397);
     when "000110001110" => data <= triangle_rom(398);
     when "000110001111" => data <= triangle_rom(399);
     when "000110010000" => data <= triangle_rom(400);
     when "000110010001" => data <= triangle_rom(401);
     when "000110010010" => data <= triangle_rom(402);
     when "000110010011" => data <= triangle_rom(403);
     when "000110010100" => data <= triangle_rom(404);
     when "000110010101" => data <= triangle_rom(405);
     when "000110010110" => data <= triangle_rom(406);
     when "000110010111" => data <= triangle_rom(407);
     when "000110011000" => data <= triangle_rom(408);
     when "000110011001" => data <= triangle_rom(409);
     when "000110011010" => data <= triangle_rom(410);
     when "000110011011" => data <= triangle_rom(411);
     when "000110011100" => data <= triangle_rom(412);
     when "000110011101" => data <= triangle_rom(413);
     when "000110011110" => data <= triangle_rom(414);
     when "000110011111" => data <= triangle_rom(415);
     when "000110100000" => data <= triangle_rom(416);
     when "000110100001" => data <= triangle_rom(417);
     when "000110100010" => data <= triangle_rom(418);
     when "000110100011" => data <= triangle_rom(419);
     when "000110100100" => data <= triangle_rom(420);
     when "000110100101" => data <= triangle_rom(421);
     when "000110100110" => data <= triangle_rom(422);
     when "000110100111" => data <= triangle_rom(423);
     when "000110101000" => data <= triangle_rom(424);
     when "000110101001" => data <= triangle_rom(425);
     when "000110101010" => data <= triangle_rom(426);
     when "000110101011" => data <= triangle_rom(427);
     when "000110101100" => data <= triangle_rom(428);
     when "000110101101" => data <= triangle_rom(429);
     when "000110101110" => data <= triangle_rom(430);
     when "000110101111" => data <= triangle_rom(431);
     when "000110110000" => data <= triangle_rom(432);
     when "000110110001" => data <= triangle_rom(433);
     when "000110110010" => data <= triangle_rom(434);
     when "000110110011" => data <= triangle_rom(435);
     when "000110110100" => data <= triangle_rom(436);
     when "000110110101" => data <= triangle_rom(437);
     when "000110110110" => data <= triangle_rom(438);
     when "000110110111" => data <= triangle_rom(439);
     when "000110111000" => data <= triangle_rom(440);
     when "000110111001" => data <= triangle_rom(441);
     when "000110111010" => data <= triangle_rom(442);
     when "000110111011" => data <= triangle_rom(443);
     when "000110111100" => data <= triangle_rom(444);
     when "000110111101" => data <= triangle_rom(445);
     when "000110111110" => data <= triangle_rom(446);
     when "000110111111" => data <= triangle_rom(447);
     when "000111000000" => data <= triangle_rom(448);
     when "000111000001" => data <= triangle_rom(449);
     when "000111000010" => data <= triangle_rom(450);
     when "000111000011" => data <= triangle_rom(451);
     when "000111000100" => data <= triangle_rom(452);
     when "000111000101" => data <= triangle_rom(453);
     when "000111000110" => data <= triangle_rom(454);
     when "000111000111" => data <= triangle_rom(455);
     when "000111001000" => data <= triangle_rom(456);
     when "000111001001" => data <= triangle_rom(457);
     when "000111001010" => data <= triangle_rom(458);
     when "000111001011" => data <= triangle_rom(459);
     when "000111001100" => data <= triangle_rom(460);
     when "000111001101" => data <= triangle_rom(461);
     when "000111001110" => data <= triangle_rom(462);
     when "000111001111" => data <= triangle_rom(463);
     when "000111010000" => data <= triangle_rom(464);
     when "000111010001" => data <= triangle_rom(465);
     when "000111010010" => data <= triangle_rom(466);
     when "000111010011" => data <= triangle_rom(467);
     when "000111010100" => data <= triangle_rom(468);
     when "000111010101" => data <= triangle_rom(469);
     when "000111010110" => data <= triangle_rom(470);
     when "000111010111" => data <= triangle_rom(471);
     when "000111011000" => data <= triangle_rom(472);
     when "000111011001" => data <= triangle_rom(473);
     when "000111011010" => data <= triangle_rom(474);
     when "000111011011" => data <= triangle_rom(475);
     when "000111011100" => data <= triangle_rom(476);
     when "000111011101" => data <= triangle_rom(477);
     when "000111011110" => data <= triangle_rom(478);
     when "000111011111" => data <= triangle_rom(479);
     when "000111100000" => data <= triangle_rom(480);
     when "000111100001" => data <= triangle_rom(481);
     when "000111100010" => data <= triangle_rom(482);
     when "000111100011" => data <= triangle_rom(483);
     when "000111100100" => data <= triangle_rom(484);
     when "000111100101" => data <= triangle_rom(485);
     when "000111100110" => data <= triangle_rom(486);
     when "000111100111" => data <= triangle_rom(487);
     when "000111101000" => data <= triangle_rom(488);
     when "000111101001" => data <= triangle_rom(489);
     when "000111101010" => data <= triangle_rom(490);
     when "000111101011" => data <= triangle_rom(491);
     when "000111101100" => data <= triangle_rom(492);
     when "000111101101" => data <= triangle_rom(493);
     when "000111101110" => data <= triangle_rom(494);
     when "000111101111" => data <= triangle_rom(495);
     when "000111110000" => data <= triangle_rom(496);
     when "000111110001" => data <= triangle_rom(497);
     when "000111110010" => data <= triangle_rom(498);
     when "000111110011" => data <= triangle_rom(499);
     when "000111110100" => data <= triangle_rom(500);
     when "000111110101" => data <= triangle_rom(501);
     when "000111110110" => data <= triangle_rom(502);
     when "000111110111" => data <= triangle_rom(503);
     when "000111111000" => data <= triangle_rom(504);
     when "000111111001" => data <= triangle_rom(505);
     when "000111111010" => data <= triangle_rom(506);
     when "000111111011" => data <= triangle_rom(507);
     when "000111111100" => data <= triangle_rom(508);
     when "000111111101" => data <= triangle_rom(509);
     when "000111111110" => data <= triangle_rom(510);
     when "000111111111" => data <= triangle_rom(511);
     when "001000000000" => data <= triangle_rom(512);
     when "001000000001" => data <= triangle_rom(513);
     when "001000000010" => data <= triangle_rom(514);
     when "001000000011" => data <= triangle_rom(515);
     when "001000000100" => data <= triangle_rom(516);
     when "001000000101" => data <= triangle_rom(517);
     when "001000000110" => data <= triangle_rom(518);
     when "001000000111" => data <= triangle_rom(519);
     when "001000001000" => data <= triangle_rom(520);
     when "001000001001" => data <= triangle_rom(521);
     when "001000001010" => data <= triangle_rom(522);
     when "001000001011" => data <= triangle_rom(523);
     when "001000001100" => data <= triangle_rom(524);
     when "001000001101" => data <= triangle_rom(525);
     when "001000001110" => data <= triangle_rom(526);
     when "001000001111" => data <= triangle_rom(527);
     when "001000010000" => data <= triangle_rom(528);
     when "001000010001" => data <= triangle_rom(529);
     when "001000010010" => data <= triangle_rom(530);
     when "001000010011" => data <= triangle_rom(531);
     when "001000010100" => data <= triangle_rom(532);
     when "001000010101" => data <= triangle_rom(533);
     when "001000010110" => data <= triangle_rom(534);
     when "001000010111" => data <= triangle_rom(535);
     when "001000011000" => data <= triangle_rom(536);
     when "001000011001" => data <= triangle_rom(537);
     when "001000011010" => data <= triangle_rom(538);
     when "001000011011" => data <= triangle_rom(539);
     when "001000011100" => data <= triangle_rom(540);
     when "001000011101" => data <= triangle_rom(541);
     when "001000011110" => data <= triangle_rom(542);
     when "001000011111" => data <= triangle_rom(543);
     when "001000100000" => data <= triangle_rom(544);
     when "001000100001" => data <= triangle_rom(545);
     when "001000100010" => data <= triangle_rom(546);
     when "001000100011" => data <= triangle_rom(547);
     when "001000100100" => data <= triangle_rom(548);
     when "001000100101" => data <= triangle_rom(549);
     when "001000100110" => data <= triangle_rom(550);
     when "001000100111" => data <= triangle_rom(551);
     when "001000101000" => data <= triangle_rom(552);
     when "001000101001" => data <= triangle_rom(553);
     when "001000101010" => data <= triangle_rom(554);
     when "001000101011" => data <= triangle_rom(555);
     when "001000101100" => data <= triangle_rom(556);
     when "001000101101" => data <= triangle_rom(557);
     when "001000101110" => data <= triangle_rom(558);
     when "001000101111" => data <= triangle_rom(559);
     when "001000110000" => data <= triangle_rom(560);
     when "001000110001" => data <= triangle_rom(561);
     when "001000110010" => data <= triangle_rom(562);
     when "001000110011" => data <= triangle_rom(563);
     when "001000110100" => data <= triangle_rom(564);
     when "001000110101" => data <= triangle_rom(565);
     when "001000110110" => data <= triangle_rom(566);
     when "001000110111" => data <= triangle_rom(567);
     when "001000111000" => data <= triangle_rom(568);
     when "001000111001" => data <= triangle_rom(569);
     when "001000111010" => data <= triangle_rom(570);
     when "001000111011" => data <= triangle_rom(571);
     when "001000111100" => data <= triangle_rom(572);
     when "001000111101" => data <= triangle_rom(573);
     when "001000111110" => data <= triangle_rom(574);
     when "001000111111" => data <= triangle_rom(575);
     when "001001000000" => data <= triangle_rom(576);
     when "001001000001" => data <= triangle_rom(577);
     when "001001000010" => data <= triangle_rom(578);
     when "001001000011" => data <= triangle_rom(579);
     when "001001000100" => data <= triangle_rom(580);
     when "001001000101" => data <= triangle_rom(581);
     when "001001000110" => data <= triangle_rom(582);
     when "001001000111" => data <= triangle_rom(583);
     when "001001001000" => data <= triangle_rom(584);
     when "001001001001" => data <= triangle_rom(585);
     when "001001001010" => data <= triangle_rom(586);
     when "001001001011" => data <= triangle_rom(587);
     when "001001001100" => data <= triangle_rom(588);
     when "001001001101" => data <= triangle_rom(589);
     when "001001001110" => data <= triangle_rom(590);
     when "001001001111" => data <= triangle_rom(591);
     when "001001010000" => data <= triangle_rom(592);
     when "001001010001" => data <= triangle_rom(593);
     when "001001010010" => data <= triangle_rom(594);
     when "001001010011" => data <= triangle_rom(595);
     when "001001010100" => data <= triangle_rom(596);
     when "001001010101" => data <= triangle_rom(597);
     when "001001010110" => data <= triangle_rom(598);
     when "001001010111" => data <= triangle_rom(599);
     when "001001011000" => data <= triangle_rom(600);
     when "001001011001" => data <= triangle_rom(601);
     when "001001011010" => data <= triangle_rom(602);
     when "001001011011" => data <= triangle_rom(603);
     when "001001011100" => data <= triangle_rom(604);
     when "001001011101" => data <= triangle_rom(605);
     when "001001011110" => data <= triangle_rom(606);
     when "001001011111" => data <= triangle_rom(607);
     when "001001100000" => data <= triangle_rom(608);
     when "001001100001" => data <= triangle_rom(609);
     when "001001100010" => data <= triangle_rom(610);
     when "001001100011" => data <= triangle_rom(611);
     when "001001100100" => data <= triangle_rom(612);
     when "001001100101" => data <= triangle_rom(613);
     when "001001100110" => data <= triangle_rom(614);
     when "001001100111" => data <= triangle_rom(615);
     when "001001101000" => data <= triangle_rom(616);
     when "001001101001" => data <= triangle_rom(617);
     when "001001101010" => data <= triangle_rom(618);
     when "001001101011" => data <= triangle_rom(619);
     when "001001101100" => data <= triangle_rom(620);
     when "001001101101" => data <= triangle_rom(621);
     when "001001101110" => data <= triangle_rom(622);
     when "001001101111" => data <= triangle_rom(623);
     when "001001110000" => data <= triangle_rom(624);
     when "001001110001" => data <= triangle_rom(625);
     when "001001110010" => data <= triangle_rom(626);
     when "001001110011" => data <= triangle_rom(627);
     when "001001110100" => data <= triangle_rom(628);
     when "001001110101" => data <= triangle_rom(629);
     when "001001110110" => data <= triangle_rom(630);
     when "001001110111" => data <= triangle_rom(631);
     when "001001111000" => data <= triangle_rom(632);
     when "001001111001" => data <= triangle_rom(633);
     when "001001111010" => data <= triangle_rom(634);
     when "001001111011" => data <= triangle_rom(635);
     when "001001111100" => data <= triangle_rom(636);
     when "001001111101" => data <= triangle_rom(637);
     when "001001111110" => data <= triangle_rom(638);
     when "001001111111" => data <= triangle_rom(639);
     when "001010000000" => data <= triangle_rom(640);
     when "001010000001" => data <= triangle_rom(641);
     when "001010000010" => data <= triangle_rom(642);
     when "001010000011" => data <= triangle_rom(643);
     when "001010000100" => data <= triangle_rom(644);
     when "001010000101" => data <= triangle_rom(645);
     when "001010000110" => data <= triangle_rom(646);
     when "001010000111" => data <= triangle_rom(647);
     when "001010001000" => data <= triangle_rom(648);
     when "001010001001" => data <= triangle_rom(649);
     when "001010001010" => data <= triangle_rom(650);
     when "001010001011" => data <= triangle_rom(651);
     when "001010001100" => data <= triangle_rom(652);
     when "001010001101" => data <= triangle_rom(653);
     when "001010001110" => data <= triangle_rom(654);
     when "001010001111" => data <= triangle_rom(655);
     when "001010010000" => data <= triangle_rom(656);
     when "001010010001" => data <= triangle_rom(657);
     when "001010010010" => data <= triangle_rom(658);
     when "001010010011" => data <= triangle_rom(659);
     when "001010010100" => data <= triangle_rom(660);
     when "001010010101" => data <= triangle_rom(661);
     when "001010010110" => data <= triangle_rom(662);
     when "001010010111" => data <= triangle_rom(663);
     when "001010011000" => data <= triangle_rom(664);
     when "001010011001" => data <= triangle_rom(665);
     when "001010011010" => data <= triangle_rom(666);
     when "001010011011" => data <= triangle_rom(667);
     when "001010011100" => data <= triangle_rom(668);
     when "001010011101" => data <= triangle_rom(669);
     when "001010011110" => data <= triangle_rom(670);
     when "001010011111" => data <= triangle_rom(671);
     when "001010100000" => data <= triangle_rom(672);
     when "001010100001" => data <= triangle_rom(673);
     when "001010100010" => data <= triangle_rom(674);
     when "001010100011" => data <= triangle_rom(675);
     when "001010100100" => data <= triangle_rom(676);
     when "001010100101" => data <= triangle_rom(677);
     when "001010100110" => data <= triangle_rom(678);
     when "001010100111" => data <= triangle_rom(679);
     when "001010101000" => data <= triangle_rom(680);
     when "001010101001" => data <= triangle_rom(681);
     when "001010101010" => data <= triangle_rom(682);
     when "001010101011" => data <= triangle_rom(683);
     when "001010101100" => data <= triangle_rom(684);
     when "001010101101" => data <= triangle_rom(685);
     when "001010101110" => data <= triangle_rom(686);
     when "001010101111" => data <= triangle_rom(687);
     when "001010110000" => data <= triangle_rom(688);
     when "001010110001" => data <= triangle_rom(689);
     when "001010110010" => data <= triangle_rom(690);
     when "001010110011" => data <= triangle_rom(691);
     when "001010110100" => data <= triangle_rom(692);
     when "001010110101" => data <= triangle_rom(693);
     when "001010110110" => data <= triangle_rom(694);
     when "001010110111" => data <= triangle_rom(695);
     when "001010111000" => data <= triangle_rom(696);
     when "001010111001" => data <= triangle_rom(697);
     when "001010111010" => data <= triangle_rom(698);
     when "001010111011" => data <= triangle_rom(699);
     when "001010111100" => data <= triangle_rom(700);
     when "001010111101" => data <= triangle_rom(701);
     when "001010111110" => data <= triangle_rom(702);
     when "001010111111" => data <= triangle_rom(703);
     when "001011000000" => data <= triangle_rom(704);
     when "001011000001" => data <= triangle_rom(705);
     when "001011000010" => data <= triangle_rom(706);
     when "001011000011" => data <= triangle_rom(707);
     when "001011000100" => data <= triangle_rom(708);
     when "001011000101" => data <= triangle_rom(709);
     when "001011000110" => data <= triangle_rom(710);
     when "001011000111" => data <= triangle_rom(711);
     when "001011001000" => data <= triangle_rom(712);
     when "001011001001" => data <= triangle_rom(713);
     when "001011001010" => data <= triangle_rom(714);
     when "001011001011" => data <= triangle_rom(715);
     when "001011001100" => data <= triangle_rom(716);
     when "001011001101" => data <= triangle_rom(717);
     when "001011001110" => data <= triangle_rom(718);
     when "001011001111" => data <= triangle_rom(719);
     when "001011010000" => data <= triangle_rom(720);
     when "001011010001" => data <= triangle_rom(721);
     when "001011010010" => data <= triangle_rom(722);
     when "001011010011" => data <= triangle_rom(723);
     when "001011010100" => data <= triangle_rom(724);
     when "001011010101" => data <= triangle_rom(725);
     when "001011010110" => data <= triangle_rom(726);
     when "001011010111" => data <= triangle_rom(727);
     when "001011011000" => data <= triangle_rom(728);
     when "001011011001" => data <= triangle_rom(729);
     when "001011011010" => data <= triangle_rom(730);
     when "001011011011" => data <= triangle_rom(731);
     when "001011011100" => data <= triangle_rom(732);
     when "001011011101" => data <= triangle_rom(733);
     when "001011011110" => data <= triangle_rom(734);
     when "001011011111" => data <= triangle_rom(735);
     when "001011100000" => data <= triangle_rom(736);
     when "001011100001" => data <= triangle_rom(737);
     when "001011100010" => data <= triangle_rom(738);
     when "001011100011" => data <= triangle_rom(739);
     when "001011100100" => data <= triangle_rom(740);
     when "001011100101" => data <= triangle_rom(741);
     when "001011100110" => data <= triangle_rom(742);
     when "001011100111" => data <= triangle_rom(743);
     when "001011101000" => data <= triangle_rom(744);
     when "001011101001" => data <= triangle_rom(745);
     when "001011101010" => data <= triangle_rom(746);
     when "001011101011" => data <= triangle_rom(747);
     when "001011101100" => data <= triangle_rom(748);
     when "001011101101" => data <= triangle_rom(749);
     when "001011101110" => data <= triangle_rom(750);
     when "001011101111" => data <= triangle_rom(751);
     when "001011110000" => data <= triangle_rom(752);
     when "001011110001" => data <= triangle_rom(753);
     when "001011110010" => data <= triangle_rom(754);
     when "001011110011" => data <= triangle_rom(755);
     when "001011110100" => data <= triangle_rom(756);
     when "001011110101" => data <= triangle_rom(757);
     when "001011110110" => data <= triangle_rom(758);
     when "001011110111" => data <= triangle_rom(759);
     when "001011111000" => data <= triangle_rom(760);
     when "001011111001" => data <= triangle_rom(761);
     when "001011111010" => data <= triangle_rom(762);
     when "001011111011" => data <= triangle_rom(763);
     when "001011111100" => data <= triangle_rom(764);
     when "001011111101" => data <= triangle_rom(765);
     when "001011111110" => data <= triangle_rom(766);
     when "001011111111" => data <= triangle_rom(767);
     when "001100000000" => data <= triangle_rom(768);
     when "001100000001" => data <= triangle_rom(769);
     when "001100000010" => data <= triangle_rom(770);
     when "001100000011" => data <= triangle_rom(771);
     when "001100000100" => data <= triangle_rom(772);
     when "001100000101" => data <= triangle_rom(773);
     when "001100000110" => data <= triangle_rom(774);
     when "001100000111" => data <= triangle_rom(775);
     when "001100001000" => data <= triangle_rom(776);
     when "001100001001" => data <= triangle_rom(777);
     when "001100001010" => data <= triangle_rom(778);
     when "001100001011" => data <= triangle_rom(779);
     when "001100001100" => data <= triangle_rom(780);
     when "001100001101" => data <= triangle_rom(781);
     when "001100001110" => data <= triangle_rom(782);
     when "001100001111" => data <= triangle_rom(783);
     when "001100010000" => data <= triangle_rom(784);
     when "001100010001" => data <= triangle_rom(785);
     when "001100010010" => data <= triangle_rom(786);
     when "001100010011" => data <= triangle_rom(787);
     when "001100010100" => data <= triangle_rom(788);
     when "001100010101" => data <= triangle_rom(789);
     when "001100010110" => data <= triangle_rom(790);
     when "001100010111" => data <= triangle_rom(791);
     when "001100011000" => data <= triangle_rom(792);
     when "001100011001" => data <= triangle_rom(793);
     when "001100011010" => data <= triangle_rom(794);
     when "001100011011" => data <= triangle_rom(795);
     when "001100011100" => data <= triangle_rom(796);
     when "001100011101" => data <= triangle_rom(797);
     when "001100011110" => data <= triangle_rom(798);
     when "001100011111" => data <= triangle_rom(799);
     when "001100100000" => data <= triangle_rom(800);
     when "001100100001" => data <= triangle_rom(801);
     when "001100100010" => data <= triangle_rom(802);
     when "001100100011" => data <= triangle_rom(803);
     when "001100100100" => data <= triangle_rom(804);
     when "001100100101" => data <= triangle_rom(805);
     when "001100100110" => data <= triangle_rom(806);
     when "001100100111" => data <= triangle_rom(807);
     when "001100101000" => data <= triangle_rom(808);
     when "001100101001" => data <= triangle_rom(809);
     when "001100101010" => data <= triangle_rom(810);
     when "001100101011" => data <= triangle_rom(811);
     when "001100101100" => data <= triangle_rom(812);
     when "001100101101" => data <= triangle_rom(813);
     when "001100101110" => data <= triangle_rom(814);
     when "001100101111" => data <= triangle_rom(815);
     when "001100110000" => data <= triangle_rom(816);
     when "001100110001" => data <= triangle_rom(817);
     when "001100110010" => data <= triangle_rom(818);
     when "001100110011" => data <= triangle_rom(819);
     when "001100110100" => data <= triangle_rom(820);
     when "001100110101" => data <= triangle_rom(821);
     when "001100110110" => data <= triangle_rom(822);
     when "001100110111" => data <= triangle_rom(823);
     when "001100111000" => data <= triangle_rom(824);
     when "001100111001" => data <= triangle_rom(825);
     when "001100111010" => data <= triangle_rom(826);
     when "001100111011" => data <= triangle_rom(827);
     when "001100111100" => data <= triangle_rom(828);
     when "001100111101" => data <= triangle_rom(829);
     when "001100111110" => data <= triangle_rom(830);
     when "001100111111" => data <= triangle_rom(831);
     when "001101000000" => data <= triangle_rom(832);
     when "001101000001" => data <= triangle_rom(833);
     when "001101000010" => data <= triangle_rom(834);
     when "001101000011" => data <= triangle_rom(835);
     when "001101000100" => data <= triangle_rom(836);
     when "001101000101" => data <= triangle_rom(837);
     when "001101000110" => data <= triangle_rom(838);
     when "001101000111" => data <= triangle_rom(839);
     when "001101001000" => data <= triangle_rom(840);
     when "001101001001" => data <= triangle_rom(841);
     when "001101001010" => data <= triangle_rom(842);
     when "001101001011" => data <= triangle_rom(843);
     when "001101001100" => data <= triangle_rom(844);
     when "001101001101" => data <= triangle_rom(845);
     when "001101001110" => data <= triangle_rom(846);
     when "001101001111" => data <= triangle_rom(847);
     when "001101010000" => data <= triangle_rom(848);
     when "001101010001" => data <= triangle_rom(849);
     when "001101010010" => data <= triangle_rom(850);
     when "001101010011" => data <= triangle_rom(851);
     when "001101010100" => data <= triangle_rom(852);
     when "001101010101" => data <= triangle_rom(853);
     when "001101010110" => data <= triangle_rom(854);
     when "001101010111" => data <= triangle_rom(855);
     when "001101011000" => data <= triangle_rom(856);
     when "001101011001" => data <= triangle_rom(857);
     when "001101011010" => data <= triangle_rom(858);
     when "001101011011" => data <= triangle_rom(859);
     when "001101011100" => data <= triangle_rom(860);
     when "001101011101" => data <= triangle_rom(861);
     when "001101011110" => data <= triangle_rom(862);
     when "001101011111" => data <= triangle_rom(863);
     when "001101100000" => data <= triangle_rom(864);
     when "001101100001" => data <= triangle_rom(865);
     when "001101100010" => data <= triangle_rom(866);
     when "001101100011" => data <= triangle_rom(867);
     when "001101100100" => data <= triangle_rom(868);
     when "001101100101" => data <= triangle_rom(869);
     when "001101100110" => data <= triangle_rom(870);
     when "001101100111" => data <= triangle_rom(871);
     when "001101101000" => data <= triangle_rom(872);
     when "001101101001" => data <= triangle_rom(873);
     when "001101101010" => data <= triangle_rom(874);
     when "001101101011" => data <= triangle_rom(875);
     when "001101101100" => data <= triangle_rom(876);
     when "001101101101" => data <= triangle_rom(877);
     when "001101101110" => data <= triangle_rom(878);
     when "001101101111" => data <= triangle_rom(879);
     when "001101110000" => data <= triangle_rom(880);
     when "001101110001" => data <= triangle_rom(881);
     when "001101110010" => data <= triangle_rom(882);
     when "001101110011" => data <= triangle_rom(883);
     when "001101110100" => data <= triangle_rom(884);
     when "001101110101" => data <= triangle_rom(885);
     when "001101110110" => data <= triangle_rom(886);
     when "001101110111" => data <= triangle_rom(887);
     when "001101111000" => data <= triangle_rom(888);
     when "001101111001" => data <= triangle_rom(889);
     when "001101111010" => data <= triangle_rom(890);
     when "001101111011" => data <= triangle_rom(891);
     when "001101111100" => data <= triangle_rom(892);
     when "001101111101" => data <= triangle_rom(893);
     when "001101111110" => data <= triangle_rom(894);
     when "001101111111" => data <= triangle_rom(895);
     when "001110000000" => data <= triangle_rom(896);
     when "001110000001" => data <= triangle_rom(897);
     when "001110000010" => data <= triangle_rom(898);
     when "001110000011" => data <= triangle_rom(899);
     when "001110000100" => data <= triangle_rom(900);
     when "001110000101" => data <= triangle_rom(901);
     when "001110000110" => data <= triangle_rom(902);
     when "001110000111" => data <= triangle_rom(903);
     when "001110001000" => data <= triangle_rom(904);
     when "001110001001" => data <= triangle_rom(905);
     when "001110001010" => data <= triangle_rom(906);
     when "001110001011" => data <= triangle_rom(907);
     when "001110001100" => data <= triangle_rom(908);
     when "001110001101" => data <= triangle_rom(909);
     when "001110001110" => data <= triangle_rom(910);
     when "001110001111" => data <= triangle_rom(911);
     when "001110010000" => data <= triangle_rom(912);
     when "001110010001" => data <= triangle_rom(913);
     when "001110010010" => data <= triangle_rom(914);
     when "001110010011" => data <= triangle_rom(915);
     when "001110010100" => data <= triangle_rom(916);
     when "001110010101" => data <= triangle_rom(917);
     when "001110010110" => data <= triangle_rom(918);
     when "001110010111" => data <= triangle_rom(919);
     when "001110011000" => data <= triangle_rom(920);
     when "001110011001" => data <= triangle_rom(921);
     when "001110011010" => data <= triangle_rom(922);
     when "001110011011" => data <= triangle_rom(923);
     when "001110011100" => data <= triangle_rom(924);
     when "001110011101" => data <= triangle_rom(925);
     when "001110011110" => data <= triangle_rom(926);
     when "001110011111" => data <= triangle_rom(927);
     when "001110100000" => data <= triangle_rom(928);
     when "001110100001" => data <= triangle_rom(929);
     when "001110100010" => data <= triangle_rom(930);
     when "001110100011" => data <= triangle_rom(931);
     when "001110100100" => data <= triangle_rom(932);
     when "001110100101" => data <= triangle_rom(933);
     when "001110100110" => data <= triangle_rom(934);
     when "001110100111" => data <= triangle_rom(935);
     when "001110101000" => data <= triangle_rom(936);
     when "001110101001" => data <= triangle_rom(937);
     when "001110101010" => data <= triangle_rom(938);
     when "001110101011" => data <= triangle_rom(939);
     when "001110101100" => data <= triangle_rom(940);
     when "001110101101" => data <= triangle_rom(941);
     when "001110101110" => data <= triangle_rom(942);
     when "001110101111" => data <= triangle_rom(943);
     when "001110110000" => data <= triangle_rom(944);
     when "001110110001" => data <= triangle_rom(945);
     when "001110110010" => data <= triangle_rom(946);
     when "001110110011" => data <= triangle_rom(947);
     when "001110110100" => data <= triangle_rom(948);
     when "001110110101" => data <= triangle_rom(949);
     when "001110110110" => data <= triangle_rom(950);
     when "001110110111" => data <= triangle_rom(951);
     when "001110111000" => data <= triangle_rom(952);
     when "001110111001" => data <= triangle_rom(953);
     when "001110111010" => data <= triangle_rom(954);
     when "001110111011" => data <= triangle_rom(955);
     when "001110111100" => data <= triangle_rom(956);
     when "001110111101" => data <= triangle_rom(957);
     when "001110111110" => data <= triangle_rom(958);
     when "001110111111" => data <= triangle_rom(959);
     when "001111000000" => data <= triangle_rom(960);
     when "001111000001" => data <= triangle_rom(961);
     when "001111000010" => data <= triangle_rom(962);
     when "001111000011" => data <= triangle_rom(963);
     when "001111000100" => data <= triangle_rom(964);
     when "001111000101" => data <= triangle_rom(965);
     when "001111000110" => data <= triangle_rom(966);
     when "001111000111" => data <= triangle_rom(967);
     when "001111001000" => data <= triangle_rom(968);
     when "001111001001" => data <= triangle_rom(969);
     when "001111001010" => data <= triangle_rom(970);
     when "001111001011" => data <= triangle_rom(971);
     when "001111001100" => data <= triangle_rom(972);
     when "001111001101" => data <= triangle_rom(973);
     when "001111001110" => data <= triangle_rom(974);
     when "001111001111" => data <= triangle_rom(975);
     when "001111010000" => data <= triangle_rom(976);
     when "001111010001" => data <= triangle_rom(977);
     when "001111010010" => data <= triangle_rom(978);
     when "001111010011" => data <= triangle_rom(979);
     when "001111010100" => data <= triangle_rom(980);
     when "001111010101" => data <= triangle_rom(981);
     when "001111010110" => data <= triangle_rom(982);
     when "001111010111" => data <= triangle_rom(983);
     when "001111011000" => data <= triangle_rom(984);
     when "001111011001" => data <= triangle_rom(985);
     when "001111011010" => data <= triangle_rom(986);
     when "001111011011" => data <= triangle_rom(987);
     when "001111011100" => data <= triangle_rom(988);
     when "001111011101" => data <= triangle_rom(989);
     when "001111011110" => data <= triangle_rom(990);
     when "001111011111" => data <= triangle_rom(991);
     when "001111100000" => data <= triangle_rom(992);
     when "001111100001" => data <= triangle_rom(993);
     when "001111100010" => data <= triangle_rom(994);
     when "001111100011" => data <= triangle_rom(995);
     when "001111100100" => data <= triangle_rom(996);
     when "001111100101" => data <= triangle_rom(997);
     when "001111100110" => data <= triangle_rom(998);
     when "001111100111" => data <= triangle_rom(999);
     when "001111101000" => data <= triangle_rom(1000);
     when "001111101001" => data <= triangle_rom(1001);
     when "001111101010" => data <= triangle_rom(1002);
     when "001111101011" => data <= triangle_rom(1003);
     when "001111101100" => data <= triangle_rom(1004);
     when "001111101101" => data <= triangle_rom(1005);
     when "001111101110" => data <= triangle_rom(1006);
     when "001111101111" => data <= triangle_rom(1007);
     when "001111110000" => data <= triangle_rom(1008);
     when "001111110001" => data <= triangle_rom(1009);
     when "001111110010" => data <= triangle_rom(1010);
     when "001111110011" => data <= triangle_rom(1011);
     when "001111110100" => data <= triangle_rom(1012);
     when "001111110101" => data <= triangle_rom(1013);
     when "001111110110" => data <= triangle_rom(1014);
     when "001111110111" => data <= triangle_rom(1015);
     when "001111111000" => data <= triangle_rom(1016);
     when "001111111001" => data <= triangle_rom(1017);
     when "001111111010" => data <= triangle_rom(1018);
     when "001111111011" => data <= triangle_rom(1019);
     when "001111111100" => data <= triangle_rom(1020);
     when "001111111101" => data <= triangle_rom(1021);
     when "001111111110" => data <= triangle_rom(1022);
     when "001111111111" => data <= triangle_rom(1023);
     when "010000000000" => data <= triangle_rom(1024);
     when "010000000001" => data <= triangle_rom(1025);
     when "010000000010" => data <= triangle_rom(1026);
     when "010000000011" => data <= triangle_rom(1027);
     when "010000000100" => data <= triangle_rom(1028);
     when "010000000101" => data <= triangle_rom(1029);
     when "010000000110" => data <= triangle_rom(1030);
     when "010000000111" => data <= triangle_rom(1031);
     when "010000001000" => data <= triangle_rom(1032);
     when "010000001001" => data <= triangle_rom(1033);
     when "010000001010" => data <= triangle_rom(1034);
     when "010000001011" => data <= triangle_rom(1035);
     when "010000001100" => data <= triangle_rom(1036);
     when "010000001101" => data <= triangle_rom(1037);
     when "010000001110" => data <= triangle_rom(1038);
     when "010000001111" => data <= triangle_rom(1039);
     when "010000010000" => data <= triangle_rom(1040);
     when "010000010001" => data <= triangle_rom(1041);
     when "010000010010" => data <= triangle_rom(1042);
     when "010000010011" => data <= triangle_rom(1043);
     when "010000010100" => data <= triangle_rom(1044);
     when "010000010101" => data <= triangle_rom(1045);
     when "010000010110" => data <= triangle_rom(1046);
     when "010000010111" => data <= triangle_rom(1047);
     when "010000011000" => data <= triangle_rom(1048);
     when "010000011001" => data <= triangle_rom(1049);
     when "010000011010" => data <= triangle_rom(1050);
     when "010000011011" => data <= triangle_rom(1051);
     when "010000011100" => data <= triangle_rom(1052);
     when "010000011101" => data <= triangle_rom(1053);
     when "010000011110" => data <= triangle_rom(1054);
     when "010000011111" => data <= triangle_rom(1055);
     when "010000100000" => data <= triangle_rom(1056);
     when "010000100001" => data <= triangle_rom(1057);
     when "010000100010" => data <= triangle_rom(1058);
     when "010000100011" => data <= triangle_rom(1059);
     when "010000100100" => data <= triangle_rom(1060);
     when "010000100101" => data <= triangle_rom(1061);
     when "010000100110" => data <= triangle_rom(1062);
     when "010000100111" => data <= triangle_rom(1063);
     when "010000101000" => data <= triangle_rom(1064);
     when "010000101001" => data <= triangle_rom(1065);
     when "010000101010" => data <= triangle_rom(1066);
     when "010000101011" => data <= triangle_rom(1067);
     when "010000101100" => data <= triangle_rom(1068);
     when "010000101101" => data <= triangle_rom(1069);
     when "010000101110" => data <= triangle_rom(1070);
     when "010000101111" => data <= triangle_rom(1071);
     when "010000110000" => data <= triangle_rom(1072);
     when "010000110001" => data <= triangle_rom(1073);
     when "010000110010" => data <= triangle_rom(1074);
     when "010000110011" => data <= triangle_rom(1075);
     when "010000110100" => data <= triangle_rom(1076);
     when "010000110101" => data <= triangle_rom(1077);
     when "010000110110" => data <= triangle_rom(1078);
     when "010000110111" => data <= triangle_rom(1079);
     when "010000111000" => data <= triangle_rom(1080);
     when "010000111001" => data <= triangle_rom(1081);
     when "010000111010" => data <= triangle_rom(1082);
     when "010000111011" => data <= triangle_rom(1083);
     when "010000111100" => data <= triangle_rom(1084);
     when "010000111101" => data <= triangle_rom(1085);
     when "010000111110" => data <= triangle_rom(1086);
     when "010000111111" => data <= triangle_rom(1087);
     when "010001000000" => data <= triangle_rom(1088);
     when "010001000001" => data <= triangle_rom(1089);
     when "010001000010" => data <= triangle_rom(1090);
     when "010001000011" => data <= triangle_rom(1091);
     when "010001000100" => data <= triangle_rom(1092);
     when "010001000101" => data <= triangle_rom(1093);
     when "010001000110" => data <= triangle_rom(1094);
     when "010001000111" => data <= triangle_rom(1095);
     when "010001001000" => data <= triangle_rom(1096);
     when "010001001001" => data <= triangle_rom(1097);
     when "010001001010" => data <= triangle_rom(1098);
     when "010001001011" => data <= triangle_rom(1099);
     when "010001001100" => data <= triangle_rom(1100);
     when "010001001101" => data <= triangle_rom(1101);
     when "010001001110" => data <= triangle_rom(1102);
     when "010001001111" => data <= triangle_rom(1103);
     when "010001010000" => data <= triangle_rom(1104);
     when "010001010001" => data <= triangle_rom(1105);
     when "010001010010" => data <= triangle_rom(1106);
     when "010001010011" => data <= triangle_rom(1107);
     when "010001010100" => data <= triangle_rom(1108);
     when "010001010101" => data <= triangle_rom(1109);
     when "010001010110" => data <= triangle_rom(1110);
     when "010001010111" => data <= triangle_rom(1111);
     when "010001011000" => data <= triangle_rom(1112);
     when "010001011001" => data <= triangle_rom(1113);
     when "010001011010" => data <= triangle_rom(1114);
     when "010001011011" => data <= triangle_rom(1115);
     when "010001011100" => data <= triangle_rom(1116);
     when "010001011101" => data <= triangle_rom(1117);
     when "010001011110" => data <= triangle_rom(1118);
     when "010001011111" => data <= triangle_rom(1119);
     when "010001100000" => data <= triangle_rom(1120);
     when "010001100001" => data <= triangle_rom(1121);
     when "010001100010" => data <= triangle_rom(1122);
     when "010001100011" => data <= triangle_rom(1123);
     when "010001100100" => data <= triangle_rom(1124);
     when "010001100101" => data <= triangle_rom(1125);
     when "010001100110" => data <= triangle_rom(1126);
     when "010001100111" => data <= triangle_rom(1127);
     when "010001101000" => data <= triangle_rom(1128);
     when "010001101001" => data <= triangle_rom(1129);
     when "010001101010" => data <= triangle_rom(1130);
     when "010001101011" => data <= triangle_rom(1131);
     when "010001101100" => data <= triangle_rom(1132);
     when "010001101101" => data <= triangle_rom(1133);
     when "010001101110" => data <= triangle_rom(1134);
     when "010001101111" => data <= triangle_rom(1135);
     when "010001110000" => data <= triangle_rom(1136);
     when "010001110001" => data <= triangle_rom(1137);
     when "010001110010" => data <= triangle_rom(1138);
     when "010001110011" => data <= triangle_rom(1139);
     when "010001110100" => data <= triangle_rom(1140);
     when "010001110101" => data <= triangle_rom(1141);
     when "010001110110" => data <= triangle_rom(1142);
     when "010001110111" => data <= triangle_rom(1143);
     when "010001111000" => data <= triangle_rom(1144);
     when "010001111001" => data <= triangle_rom(1145);
     when "010001111010" => data <= triangle_rom(1146);
     when "010001111011" => data <= triangle_rom(1147);
     when "010001111100" => data <= triangle_rom(1148);
     when "010001111101" => data <= triangle_rom(1149);
     when "010001111110" => data <= triangle_rom(1150);
     when "010001111111" => data <= triangle_rom(1151);
     when "010010000000" => data <= triangle_rom(1152);
     when "010010000001" => data <= triangle_rom(1153);
     when "010010000010" => data <= triangle_rom(1154);
     when "010010000011" => data <= triangle_rom(1155);
     when "010010000100" => data <= triangle_rom(1156);
     when "010010000101" => data <= triangle_rom(1157);
     when "010010000110" => data <= triangle_rom(1158);
     when "010010000111" => data <= triangle_rom(1159);
     when "010010001000" => data <= triangle_rom(1160);
     when "010010001001" => data <= triangle_rom(1161);
     when "010010001010" => data <= triangle_rom(1162);
     when "010010001011" => data <= triangle_rom(1163);
     when "010010001100" => data <= triangle_rom(1164);
     when "010010001101" => data <= triangle_rom(1165);
     when "010010001110" => data <= triangle_rom(1166);
     when "010010001111" => data <= triangle_rom(1167);
     when "010010010000" => data <= triangle_rom(1168);
     when "010010010001" => data <= triangle_rom(1169);
     when "010010010010" => data <= triangle_rom(1170);
     when "010010010011" => data <= triangle_rom(1171);
     when "010010010100" => data <= triangle_rom(1172);
     when "010010010101" => data <= triangle_rom(1173);
     when "010010010110" => data <= triangle_rom(1174);
     when "010010010111" => data <= triangle_rom(1175);
     when "010010011000" => data <= triangle_rom(1176);
     when "010010011001" => data <= triangle_rom(1177);
     when "010010011010" => data <= triangle_rom(1178);
     when "010010011011" => data <= triangle_rom(1179);
     when "010010011100" => data <= triangle_rom(1180);
     when "010010011101" => data <= triangle_rom(1181);
     when "010010011110" => data <= triangle_rom(1182);
     when "010010011111" => data <= triangle_rom(1183);
     when "010010100000" => data <= triangle_rom(1184);
     when "010010100001" => data <= triangle_rom(1185);
     when "010010100010" => data <= triangle_rom(1186);
     when "010010100011" => data <= triangle_rom(1187);
     when "010010100100" => data <= triangle_rom(1188);
     when "010010100101" => data <= triangle_rom(1189);
     when "010010100110" => data <= triangle_rom(1190);
     when "010010100111" => data <= triangle_rom(1191);
     when "010010101000" => data <= triangle_rom(1192);
     when "010010101001" => data <= triangle_rom(1193);
     when "010010101010" => data <= triangle_rom(1194);
     when "010010101011" => data <= triangle_rom(1195);
     when "010010101100" => data <= triangle_rom(1196);
     when "010010101101" => data <= triangle_rom(1197);
     when "010010101110" => data <= triangle_rom(1198);
     when "010010101111" => data <= triangle_rom(1199);
     when "010010110000" => data <= triangle_rom(1200);
     when "010010110001" => data <= triangle_rom(1201);
     when "010010110010" => data <= triangle_rom(1202);
     when "010010110011" => data <= triangle_rom(1203);
     when "010010110100" => data <= triangle_rom(1204);
     when "010010110101" => data <= triangle_rom(1205);
     when "010010110110" => data <= triangle_rom(1206);
     when "010010110111" => data <= triangle_rom(1207);
     when "010010111000" => data <= triangle_rom(1208);
     when "010010111001" => data <= triangle_rom(1209);
     when "010010111010" => data <= triangle_rom(1210);
     when "010010111011" => data <= triangle_rom(1211);
     when "010010111100" => data <= triangle_rom(1212);
     when "010010111101" => data <= triangle_rom(1213);
     when "010010111110" => data <= triangle_rom(1214);
     when "010010111111" => data <= triangle_rom(1215);
     when "010011000000" => data <= triangle_rom(1216);
     when "010011000001" => data <= triangle_rom(1217);
     when "010011000010" => data <= triangle_rom(1218);
     when "010011000011" => data <= triangle_rom(1219);
     when "010011000100" => data <= triangle_rom(1220);
     when "010011000101" => data <= triangle_rom(1221);
     when "010011000110" => data <= triangle_rom(1222);
     when "010011000111" => data <= triangle_rom(1223);
     when "010011001000" => data <= triangle_rom(1224);
     when "010011001001" => data <= triangle_rom(1225);
     when "010011001010" => data <= triangle_rom(1226);
     when "010011001011" => data <= triangle_rom(1227);
     when "010011001100" => data <= triangle_rom(1228);
     when "010011001101" => data <= triangle_rom(1229);
     when "010011001110" => data <= triangle_rom(1230);
     when "010011001111" => data <= triangle_rom(1231);
     when "010011010000" => data <= triangle_rom(1232);
     when "010011010001" => data <= triangle_rom(1233);
     when "010011010010" => data <= triangle_rom(1234);
     when "010011010011" => data <= triangle_rom(1235);
     when "010011010100" => data <= triangle_rom(1236);
     when "010011010101" => data <= triangle_rom(1237);
     when "010011010110" => data <= triangle_rom(1238);
     when "010011010111" => data <= triangle_rom(1239);
     when "010011011000" => data <= triangle_rom(1240);
     when "010011011001" => data <= triangle_rom(1241);
     when "010011011010" => data <= triangle_rom(1242);
     when "010011011011" => data <= triangle_rom(1243);
     when "010011011100" => data <= triangle_rom(1244);
     when "010011011101" => data <= triangle_rom(1245);
     when "010011011110" => data <= triangle_rom(1246);
     when "010011011111" => data <= triangle_rom(1247);
     when "010011100000" => data <= triangle_rom(1248);
     when "010011100001" => data <= triangle_rom(1249);
     when "010011100010" => data <= triangle_rom(1250);
     when "010011100011" => data <= triangle_rom(1251);
     when "010011100100" => data <= triangle_rom(1252);
     when "010011100101" => data <= triangle_rom(1253);
     when "010011100110" => data <= triangle_rom(1254);
     when "010011100111" => data <= triangle_rom(1255);
     when "010011101000" => data <= triangle_rom(1256);
     when "010011101001" => data <= triangle_rom(1257);
     when "010011101010" => data <= triangle_rom(1258);
     when "010011101011" => data <= triangle_rom(1259);
     when "010011101100" => data <= triangle_rom(1260);
     when "010011101101" => data <= triangle_rom(1261);
     when "010011101110" => data <= triangle_rom(1262);
     when "010011101111" => data <= triangle_rom(1263);
     when "010011110000" => data <= triangle_rom(1264);
     when "010011110001" => data <= triangle_rom(1265);
     when "010011110010" => data <= triangle_rom(1266);
     when "010011110011" => data <= triangle_rom(1267);
     when "010011110100" => data <= triangle_rom(1268);
     when "010011110101" => data <= triangle_rom(1269);
     when "010011110110" => data <= triangle_rom(1270);
     when "010011110111" => data <= triangle_rom(1271);
     when "010011111000" => data <= triangle_rom(1272);
     when "010011111001" => data <= triangle_rom(1273);
     when "010011111010" => data <= triangle_rom(1274);
     when "010011111011" => data <= triangle_rom(1275);
     when "010011111100" => data <= triangle_rom(1276);
     when "010011111101" => data <= triangle_rom(1277);
     when "010011111110" => data <= triangle_rom(1278);
     when "010011111111" => data <= triangle_rom(1279);
     when "010100000000" => data <= triangle_rom(1280);
     when "010100000001" => data <= triangle_rom(1281);
     when "010100000010" => data <= triangle_rom(1282);
     when "010100000011" => data <= triangle_rom(1283);
     when "010100000100" => data <= triangle_rom(1284);
     when "010100000101" => data <= triangle_rom(1285);
     when "010100000110" => data <= triangle_rom(1286);
     when "010100000111" => data <= triangle_rom(1287);
     when "010100001000" => data <= triangle_rom(1288);
     when "010100001001" => data <= triangle_rom(1289);
     when "010100001010" => data <= triangle_rom(1290);
     when "010100001011" => data <= triangle_rom(1291);
     when "010100001100" => data <= triangle_rom(1292);
     when "010100001101" => data <= triangle_rom(1293);
     when "010100001110" => data <= triangle_rom(1294);
     when "010100001111" => data <= triangle_rom(1295);
     when "010100010000" => data <= triangle_rom(1296);
     when "010100010001" => data <= triangle_rom(1297);
     when "010100010010" => data <= triangle_rom(1298);
     when "010100010011" => data <= triangle_rom(1299);
     when "010100010100" => data <= triangle_rom(1300);
     when "010100010101" => data <= triangle_rom(1301);
     when "010100010110" => data <= triangle_rom(1302);
     when "010100010111" => data <= triangle_rom(1303);
     when "010100011000" => data <= triangle_rom(1304);
     when "010100011001" => data <= triangle_rom(1305);
     when "010100011010" => data <= triangle_rom(1306);
     when "010100011011" => data <= triangle_rom(1307);
     when "010100011100" => data <= triangle_rom(1308);
     when "010100011101" => data <= triangle_rom(1309);
     when "010100011110" => data <= triangle_rom(1310);
     when "010100011111" => data <= triangle_rom(1311);
     when "010100100000" => data <= triangle_rom(1312);
     when "010100100001" => data <= triangle_rom(1313);
     when "010100100010" => data <= triangle_rom(1314);
     when "010100100011" => data <= triangle_rom(1315);
     when "010100100100" => data <= triangle_rom(1316);
     when "010100100101" => data <= triangle_rom(1317);
     when "010100100110" => data <= triangle_rom(1318);
     when "010100100111" => data <= triangle_rom(1319);
     when "010100101000" => data <= triangle_rom(1320);
     when "010100101001" => data <= triangle_rom(1321);
     when "010100101010" => data <= triangle_rom(1322);
     when "010100101011" => data <= triangle_rom(1323);
     when "010100101100" => data <= triangle_rom(1324);
     when "010100101101" => data <= triangle_rom(1325);
     when "010100101110" => data <= triangle_rom(1326);
     when "010100101111" => data <= triangle_rom(1327);
     when "010100110000" => data <= triangle_rom(1328);
     when "010100110001" => data <= triangle_rom(1329);
     when "010100110010" => data <= triangle_rom(1330);
     when "010100110011" => data <= triangle_rom(1331);
     when "010100110100" => data <= triangle_rom(1332);
     when "010100110101" => data <= triangle_rom(1333);
     when "010100110110" => data <= triangle_rom(1334);
     when "010100110111" => data <= triangle_rom(1335);
     when "010100111000" => data <= triangle_rom(1336);
     when "010100111001" => data <= triangle_rom(1337);
     when "010100111010" => data <= triangle_rom(1338);
     when "010100111011" => data <= triangle_rom(1339);
     when "010100111100" => data <= triangle_rom(1340);
     when "010100111101" => data <= triangle_rom(1341);
     when "010100111110" => data <= triangle_rom(1342);
     when "010100111111" => data <= triangle_rom(1343);
     when "010101000000" => data <= triangle_rom(1344);
     when "010101000001" => data <= triangle_rom(1345);
     when "010101000010" => data <= triangle_rom(1346);
     when "010101000011" => data <= triangle_rom(1347);
     when "010101000100" => data <= triangle_rom(1348);
     when "010101000101" => data <= triangle_rom(1349);
     when "010101000110" => data <= triangle_rom(1350);
     when "010101000111" => data <= triangle_rom(1351);
     when "010101001000" => data <= triangle_rom(1352);
     when "010101001001" => data <= triangle_rom(1353);
     when "010101001010" => data <= triangle_rom(1354);
     when "010101001011" => data <= triangle_rom(1355);
     when "010101001100" => data <= triangle_rom(1356);
     when "010101001101" => data <= triangle_rom(1357);
     when "010101001110" => data <= triangle_rom(1358);
     when "010101001111" => data <= triangle_rom(1359);
     when "010101010000" => data <= triangle_rom(1360);
     when "010101010001" => data <= triangle_rom(1361);
     when "010101010010" => data <= triangle_rom(1362);
     when "010101010011" => data <= triangle_rom(1363);
     when "010101010100" => data <= triangle_rom(1364);
     when "010101010101" => data <= triangle_rom(1365);
     when "010101010110" => data <= triangle_rom(1366);
     when "010101010111" => data <= triangle_rom(1367);
     when "010101011000" => data <= triangle_rom(1368);
     when "010101011001" => data <= triangle_rom(1369);
     when "010101011010" => data <= triangle_rom(1370);
     when "010101011011" => data <= triangle_rom(1371);
     when "010101011100" => data <= triangle_rom(1372);
     when "010101011101" => data <= triangle_rom(1373);
     when "010101011110" => data <= triangle_rom(1374);
     when "010101011111" => data <= triangle_rom(1375);
     when "010101100000" => data <= triangle_rom(1376);
     when "010101100001" => data <= triangle_rom(1377);
     when "010101100010" => data <= triangle_rom(1378);
     when "010101100011" => data <= triangle_rom(1379);
     when "010101100100" => data <= triangle_rom(1380);
     when "010101100101" => data <= triangle_rom(1381);
     when "010101100110" => data <= triangle_rom(1382);
     when "010101100111" => data <= triangle_rom(1383);
     when "010101101000" => data <= triangle_rom(1384);
     when "010101101001" => data <= triangle_rom(1385);
     when "010101101010" => data <= triangle_rom(1386);
     when "010101101011" => data <= triangle_rom(1387);
     when "010101101100" => data <= triangle_rom(1388);
     when "010101101101" => data <= triangle_rom(1389);
     when "010101101110" => data <= triangle_rom(1390);
     when "010101101111" => data <= triangle_rom(1391);
     when "010101110000" => data <= triangle_rom(1392);
     when "010101110001" => data <= triangle_rom(1393);
     when "010101110010" => data <= triangle_rom(1394);
     when "010101110011" => data <= triangle_rom(1395);
     when "010101110100" => data <= triangle_rom(1396);
     when "010101110101" => data <= triangle_rom(1397);
     when "010101110110" => data <= triangle_rom(1398);
     when "010101110111" => data <= triangle_rom(1399);
     when "010101111000" => data <= triangle_rom(1400);
     when "010101111001" => data <= triangle_rom(1401);
     when "010101111010" => data <= triangle_rom(1402);
     when "010101111011" => data <= triangle_rom(1403);
     when "010101111100" => data <= triangle_rom(1404);
     when "010101111101" => data <= triangle_rom(1405);
     when "010101111110" => data <= triangle_rom(1406);
     when "010101111111" => data <= triangle_rom(1407);
     when "010110000000" => data <= triangle_rom(1408);
     when "010110000001" => data <= triangle_rom(1409);
     when "010110000010" => data <= triangle_rom(1410);
     when "010110000011" => data <= triangle_rom(1411);
     when "010110000100" => data <= triangle_rom(1412);
     when "010110000101" => data <= triangle_rom(1413);
     when "010110000110" => data <= triangle_rom(1414);
     when "010110000111" => data <= triangle_rom(1415);
     when "010110001000" => data <= triangle_rom(1416);
     when "010110001001" => data <= triangle_rom(1417);
     when "010110001010" => data <= triangle_rom(1418);
     when "010110001011" => data <= triangle_rom(1419);
     when "010110001100" => data <= triangle_rom(1420);
     when "010110001101" => data <= triangle_rom(1421);
     when "010110001110" => data <= triangle_rom(1422);
     when "010110001111" => data <= triangle_rom(1423);
     when "010110010000" => data <= triangle_rom(1424);
     when "010110010001" => data <= triangle_rom(1425);
     when "010110010010" => data <= triangle_rom(1426);
     when "010110010011" => data <= triangle_rom(1427);
     when "010110010100" => data <= triangle_rom(1428);
     when "010110010101" => data <= triangle_rom(1429);
     when "010110010110" => data <= triangle_rom(1430);
     when "010110010111" => data <= triangle_rom(1431);
     when "010110011000" => data <= triangle_rom(1432);
     when "010110011001" => data <= triangle_rom(1433);
     when "010110011010" => data <= triangle_rom(1434);
     when "010110011011" => data <= triangle_rom(1435);
     when "010110011100" => data <= triangle_rom(1436);
     when "010110011101" => data <= triangle_rom(1437);
     when "010110011110" => data <= triangle_rom(1438);
     when "010110011111" => data <= triangle_rom(1439);
     when "010110100000" => data <= triangle_rom(1440);
     when "010110100001" => data <= triangle_rom(1441);
     when "010110100010" => data <= triangle_rom(1442);
     when "010110100011" => data <= triangle_rom(1443);
     when "010110100100" => data <= triangle_rom(1444);
     when "010110100101" => data <= triangle_rom(1445);
     when "010110100110" => data <= triangle_rom(1446);
     when "010110100111" => data <= triangle_rom(1447);
     when "010110101000" => data <= triangle_rom(1448);
     when "010110101001" => data <= triangle_rom(1449);
     when "010110101010" => data <= triangle_rom(1450);
     when "010110101011" => data <= triangle_rom(1451);
     when "010110101100" => data <= triangle_rom(1452);
     when "010110101101" => data <= triangle_rom(1453);
     when "010110101110" => data <= triangle_rom(1454);
     when "010110101111" => data <= triangle_rom(1455);
     when "010110110000" => data <= triangle_rom(1456);
     when "010110110001" => data <= triangle_rom(1457);
     when "010110110010" => data <= triangle_rom(1458);
     when "010110110011" => data <= triangle_rom(1459);
     when "010110110100" => data <= triangle_rom(1460);
     when "010110110101" => data <= triangle_rom(1461);
     when "010110110110" => data <= triangle_rom(1462);
     when "010110110111" => data <= triangle_rom(1463);
     when "010110111000" => data <= triangle_rom(1464);
     when "010110111001" => data <= triangle_rom(1465);
     when "010110111010" => data <= triangle_rom(1466);
     when "010110111011" => data <= triangle_rom(1467);
     when "010110111100" => data <= triangle_rom(1468);
     when "010110111101" => data <= triangle_rom(1469);
     when "010110111110" => data <= triangle_rom(1470);
     when "010110111111" => data <= triangle_rom(1471);
     when "010111000000" => data <= triangle_rom(1472);
     when "010111000001" => data <= triangle_rom(1473);
     when "010111000010" => data <= triangle_rom(1474);
     when "010111000011" => data <= triangle_rom(1475);
     when "010111000100" => data <= triangle_rom(1476);
     when "010111000101" => data <= triangle_rom(1477);
     when "010111000110" => data <= triangle_rom(1478);
     when "010111000111" => data <= triangle_rom(1479);
     when "010111001000" => data <= triangle_rom(1480);
     when "010111001001" => data <= triangle_rom(1481);
     when "010111001010" => data <= triangle_rom(1482);
     when "010111001011" => data <= triangle_rom(1483);
     when "010111001100" => data <= triangle_rom(1484);
     when "010111001101" => data <= triangle_rom(1485);
     when "010111001110" => data <= triangle_rom(1486);
     when "010111001111" => data <= triangle_rom(1487);
     when "010111010000" => data <= triangle_rom(1488);
     when "010111010001" => data <= triangle_rom(1489);
     when "010111010010" => data <= triangle_rom(1490);
     when "010111010011" => data <= triangle_rom(1491);
     when "010111010100" => data <= triangle_rom(1492);
     when "010111010101" => data <= triangle_rom(1493);
     when "010111010110" => data <= triangle_rom(1494);
     when "010111010111" => data <= triangle_rom(1495);
     when "010111011000" => data <= triangle_rom(1496);
     when "010111011001" => data <= triangle_rom(1497);
     when "010111011010" => data <= triangle_rom(1498);
     when "010111011011" => data <= triangle_rom(1499);
     when "010111011100" => data <= triangle_rom(1500);
     when "010111011101" => data <= triangle_rom(1501);
     when "010111011110" => data <= triangle_rom(1502);
     when "010111011111" => data <= triangle_rom(1503);
     when "010111100000" => data <= triangle_rom(1504);
     when "010111100001" => data <= triangle_rom(1505);
     when "010111100010" => data <= triangle_rom(1506);
     when "010111100011" => data <= triangle_rom(1507);
     when "010111100100" => data <= triangle_rom(1508);
     when "010111100101" => data <= triangle_rom(1509);
     when "010111100110" => data <= triangle_rom(1510);
     when "010111100111" => data <= triangle_rom(1511);
     when "010111101000" => data <= triangle_rom(1512);
     when "010111101001" => data <= triangle_rom(1513);
     when "010111101010" => data <= triangle_rom(1514);
     when "010111101011" => data <= triangle_rom(1515);
     when "010111101100" => data <= triangle_rom(1516);
     when "010111101101" => data <= triangle_rom(1517);
     when "010111101110" => data <= triangle_rom(1518);
     when "010111101111" => data <= triangle_rom(1519);
     when "010111110000" => data <= triangle_rom(1520);
     when "010111110001" => data <= triangle_rom(1521);
     when "010111110010" => data <= triangle_rom(1522);
     when "010111110011" => data <= triangle_rom(1523);
     when "010111110100" => data <= triangle_rom(1524);
     when "010111110101" => data <= triangle_rom(1525);
     when "010111110110" => data <= triangle_rom(1526);
     when "010111110111" => data <= triangle_rom(1527);
     when "010111111000" => data <= triangle_rom(1528);
     when "010111111001" => data <= triangle_rom(1529);
     when "010111111010" => data <= triangle_rom(1530);
     when "010111111011" => data <= triangle_rom(1531);
     when "010111111100" => data <= triangle_rom(1532);
     when "010111111101" => data <= triangle_rom(1533);
     when "010111111110" => data <= triangle_rom(1534);
     when "010111111111" => data <= triangle_rom(1535);
     when "011000000000" => data <= triangle_rom(1536);
     when "011000000001" => data <= triangle_rom(1537);
     when "011000000010" => data <= triangle_rom(1538);
     when "011000000011" => data <= triangle_rom(1539);
     when "011000000100" => data <= triangle_rom(1540);
     when "011000000101" => data <= triangle_rom(1541);
     when "011000000110" => data <= triangle_rom(1542);
     when "011000000111" => data <= triangle_rom(1543);
     when "011000001000" => data <= triangle_rom(1544);
     when "011000001001" => data <= triangle_rom(1545);
     when "011000001010" => data <= triangle_rom(1546);
     when "011000001011" => data <= triangle_rom(1547);
     when "011000001100" => data <= triangle_rom(1548);
     when "011000001101" => data <= triangle_rom(1549);
     when "011000001110" => data <= triangle_rom(1550);
     when "011000001111" => data <= triangle_rom(1551);
     when "011000010000" => data <= triangle_rom(1552);
     when "011000010001" => data <= triangle_rom(1553);
     when "011000010010" => data <= triangle_rom(1554);
     when "011000010011" => data <= triangle_rom(1555);
     when "011000010100" => data <= triangle_rom(1556);
     when "011000010101" => data <= triangle_rom(1557);
     when "011000010110" => data <= triangle_rom(1558);
     when "011000010111" => data <= triangle_rom(1559);
     when "011000011000" => data <= triangle_rom(1560);
     when "011000011001" => data <= triangle_rom(1561);
     when "011000011010" => data <= triangle_rom(1562);
     when "011000011011" => data <= triangle_rom(1563);
     when "011000011100" => data <= triangle_rom(1564);
     when "011000011101" => data <= triangle_rom(1565);
     when "011000011110" => data <= triangle_rom(1566);
     when "011000011111" => data <= triangle_rom(1567);
     when "011000100000" => data <= triangle_rom(1568);
     when "011000100001" => data <= triangle_rom(1569);
     when "011000100010" => data <= triangle_rom(1570);
     when "011000100011" => data <= triangle_rom(1571);
     when "011000100100" => data <= triangle_rom(1572);
     when "011000100101" => data <= triangle_rom(1573);
     when "011000100110" => data <= triangle_rom(1574);
     when "011000100111" => data <= triangle_rom(1575);
     when "011000101000" => data <= triangle_rom(1576);
     when "011000101001" => data <= triangle_rom(1577);
     when "011000101010" => data <= triangle_rom(1578);
     when "011000101011" => data <= triangle_rom(1579);
     when "011000101100" => data <= triangle_rom(1580);
     when "011000101101" => data <= triangle_rom(1581);
     when "011000101110" => data <= triangle_rom(1582);
     when "011000101111" => data <= triangle_rom(1583);
     when "011000110000" => data <= triangle_rom(1584);
     when "011000110001" => data <= triangle_rom(1585);
     when "011000110010" => data <= triangle_rom(1586);
     when "011000110011" => data <= triangle_rom(1587);
     when "011000110100" => data <= triangle_rom(1588);
     when "011000110101" => data <= triangle_rom(1589);
     when "011000110110" => data <= triangle_rom(1590);
     when "011000110111" => data <= triangle_rom(1591);
     when "011000111000" => data <= triangle_rom(1592);
     when "011000111001" => data <= triangle_rom(1593);
     when "011000111010" => data <= triangle_rom(1594);
     when "011000111011" => data <= triangle_rom(1595);
     when "011000111100" => data <= triangle_rom(1596);
     when "011000111101" => data <= triangle_rom(1597);
     when "011000111110" => data <= triangle_rom(1598);
     when "011000111111" => data <= triangle_rom(1599);
     when "011001000000" => data <= triangle_rom(1600);
     when "011001000001" => data <= triangle_rom(1601);
     when "011001000010" => data <= triangle_rom(1602);
     when "011001000011" => data <= triangle_rom(1603);
     when "011001000100" => data <= triangle_rom(1604);
     when "011001000101" => data <= triangle_rom(1605);
     when "011001000110" => data <= triangle_rom(1606);
     when "011001000111" => data <= triangle_rom(1607);
     when "011001001000" => data <= triangle_rom(1608);
     when "011001001001" => data <= triangle_rom(1609);
     when "011001001010" => data <= triangle_rom(1610);
     when "011001001011" => data <= triangle_rom(1611);
     when "011001001100" => data <= triangle_rom(1612);
     when "011001001101" => data <= triangle_rom(1613);
     when "011001001110" => data <= triangle_rom(1614);
     when "011001001111" => data <= triangle_rom(1615);
     when "011001010000" => data <= triangle_rom(1616);
     when "011001010001" => data <= triangle_rom(1617);
     when "011001010010" => data <= triangle_rom(1618);
     when "011001010011" => data <= triangle_rom(1619);
     when "011001010100" => data <= triangle_rom(1620);
     when "011001010101" => data <= triangle_rom(1621);
     when "011001010110" => data <= triangle_rom(1622);
     when "011001010111" => data <= triangle_rom(1623);
     when "011001011000" => data <= triangle_rom(1624);
     when "011001011001" => data <= triangle_rom(1625);
     when "011001011010" => data <= triangle_rom(1626);
     when "011001011011" => data <= triangle_rom(1627);
     when "011001011100" => data <= triangle_rom(1628);
     when "011001011101" => data <= triangle_rom(1629);
     when "011001011110" => data <= triangle_rom(1630);
     when "011001011111" => data <= triangle_rom(1631);
     when "011001100000" => data <= triangle_rom(1632);
     when "011001100001" => data <= triangle_rom(1633);
     when "011001100010" => data <= triangle_rom(1634);
     when "011001100011" => data <= triangle_rom(1635);
     when "011001100100" => data <= triangle_rom(1636);
     when "011001100101" => data <= triangle_rom(1637);
     when "011001100110" => data <= triangle_rom(1638);
     when "011001100111" => data <= triangle_rom(1639);
     when "011001101000" => data <= triangle_rom(1640);
     when "011001101001" => data <= triangle_rom(1641);
     when "011001101010" => data <= triangle_rom(1642);
     when "011001101011" => data <= triangle_rom(1643);
     when "011001101100" => data <= triangle_rom(1644);
     when "011001101101" => data <= triangle_rom(1645);
     when "011001101110" => data <= triangle_rom(1646);
     when "011001101111" => data <= triangle_rom(1647);
     when "011001110000" => data <= triangle_rom(1648);
     when "011001110001" => data <= triangle_rom(1649);
     when "011001110010" => data <= triangle_rom(1650);
     when "011001110011" => data <= triangle_rom(1651);
     when "011001110100" => data <= triangle_rom(1652);
     when "011001110101" => data <= triangle_rom(1653);
     when "011001110110" => data <= triangle_rom(1654);
     when "011001110111" => data <= triangle_rom(1655);
     when "011001111000" => data <= triangle_rom(1656);
     when "011001111001" => data <= triangle_rom(1657);
     when "011001111010" => data <= triangle_rom(1658);
     when "011001111011" => data <= triangle_rom(1659);
     when "011001111100" => data <= triangle_rom(1660);
     when "011001111101" => data <= triangle_rom(1661);
     when "011001111110" => data <= triangle_rom(1662);
     when "011001111111" => data <= triangle_rom(1663);
     when "011010000000" => data <= triangle_rom(1664);
     when "011010000001" => data <= triangle_rom(1665);
     when "011010000010" => data <= triangle_rom(1666);
     when "011010000011" => data <= triangle_rom(1667);
     when "011010000100" => data <= triangle_rom(1668);
     when "011010000101" => data <= triangle_rom(1669);
     when "011010000110" => data <= triangle_rom(1670);
     when "011010000111" => data <= triangle_rom(1671);
     when "011010001000" => data <= triangle_rom(1672);
     when "011010001001" => data <= triangle_rom(1673);
     when "011010001010" => data <= triangle_rom(1674);
     when "011010001011" => data <= triangle_rom(1675);
     when "011010001100" => data <= triangle_rom(1676);
     when "011010001101" => data <= triangle_rom(1677);
     when "011010001110" => data <= triangle_rom(1678);
     when "011010001111" => data <= triangle_rom(1679);
     when "011010010000" => data <= triangle_rom(1680);
     when "011010010001" => data <= triangle_rom(1681);
     when "011010010010" => data <= triangle_rom(1682);
     when "011010010011" => data <= triangle_rom(1683);
     when "011010010100" => data <= triangle_rom(1684);
     when "011010010101" => data <= triangle_rom(1685);
     when "011010010110" => data <= triangle_rom(1686);
     when "011010010111" => data <= triangle_rom(1687);
     when "011010011000" => data <= triangle_rom(1688);
     when "011010011001" => data <= triangle_rom(1689);
     when "011010011010" => data <= triangle_rom(1690);
     when "011010011011" => data <= triangle_rom(1691);
     when "011010011100" => data <= triangle_rom(1692);
     when "011010011101" => data <= triangle_rom(1693);
     when "011010011110" => data <= triangle_rom(1694);
     when "011010011111" => data <= triangle_rom(1695);
     when "011010100000" => data <= triangle_rom(1696);
     when "011010100001" => data <= triangle_rom(1697);
     when "011010100010" => data <= triangle_rom(1698);
     when "011010100011" => data <= triangle_rom(1699);
     when "011010100100" => data <= triangle_rom(1700);
     when "011010100101" => data <= triangle_rom(1701);
     when "011010100110" => data <= triangle_rom(1702);
     when "011010100111" => data <= triangle_rom(1703);
     when "011010101000" => data <= triangle_rom(1704);
     when "011010101001" => data <= triangle_rom(1705);
     when "011010101010" => data <= triangle_rom(1706);
     when "011010101011" => data <= triangle_rom(1707);
     when "011010101100" => data <= triangle_rom(1708);
     when "011010101101" => data <= triangle_rom(1709);
     when "011010101110" => data <= triangle_rom(1710);
     when "011010101111" => data <= triangle_rom(1711);
     when "011010110000" => data <= triangle_rom(1712);
     when "011010110001" => data <= triangle_rom(1713);
     when "011010110010" => data <= triangle_rom(1714);
     when "011010110011" => data <= triangle_rom(1715);
     when "011010110100" => data <= triangle_rom(1716);
     when "011010110101" => data <= triangle_rom(1717);
     when "011010110110" => data <= triangle_rom(1718);
     when "011010110111" => data <= triangle_rom(1719);
     when "011010111000" => data <= triangle_rom(1720);
     when "011010111001" => data <= triangle_rom(1721);
     when "011010111010" => data <= triangle_rom(1722);
     when "011010111011" => data <= triangle_rom(1723);
     when "011010111100" => data <= triangle_rom(1724);
     when "011010111101" => data <= triangle_rom(1725);
     when "011010111110" => data <= triangle_rom(1726);
     when "011010111111" => data <= triangle_rom(1727);
     when "011011000000" => data <= triangle_rom(1728);
     when "011011000001" => data <= triangle_rom(1729);
     when "011011000010" => data <= triangle_rom(1730);
     when "011011000011" => data <= triangle_rom(1731);
     when "011011000100" => data <= triangle_rom(1732);
     when "011011000101" => data <= triangle_rom(1733);
     when "011011000110" => data <= triangle_rom(1734);
     when "011011000111" => data <= triangle_rom(1735);
     when "011011001000" => data <= triangle_rom(1736);
     when "011011001001" => data <= triangle_rom(1737);
     when "011011001010" => data <= triangle_rom(1738);
     when "011011001011" => data <= triangle_rom(1739);
     when "011011001100" => data <= triangle_rom(1740);
     when "011011001101" => data <= triangle_rom(1741);
     when "011011001110" => data <= triangle_rom(1742);
     when "011011001111" => data <= triangle_rom(1743);
     when "011011010000" => data <= triangle_rom(1744);
     when "011011010001" => data <= triangle_rom(1745);
     when "011011010010" => data <= triangle_rom(1746);
     when "011011010011" => data <= triangle_rom(1747);
     when "011011010100" => data <= triangle_rom(1748);
     when "011011010101" => data <= triangle_rom(1749);
     when "011011010110" => data <= triangle_rom(1750);
     when "011011010111" => data <= triangle_rom(1751);
     when "011011011000" => data <= triangle_rom(1752);
     when "011011011001" => data <= triangle_rom(1753);
     when "011011011010" => data <= triangle_rom(1754);
     when "011011011011" => data <= triangle_rom(1755);
     when "011011011100" => data <= triangle_rom(1756);
     when "011011011101" => data <= triangle_rom(1757);
     when "011011011110" => data <= triangle_rom(1758);
     when "011011011111" => data <= triangle_rom(1759);
     when "011011100000" => data <= triangle_rom(1760);
     when "011011100001" => data <= triangle_rom(1761);
     when "011011100010" => data <= triangle_rom(1762);
     when "011011100011" => data <= triangle_rom(1763);
     when "011011100100" => data <= triangle_rom(1764);
     when "011011100101" => data <= triangle_rom(1765);
     when "011011100110" => data <= triangle_rom(1766);
     when "011011100111" => data <= triangle_rom(1767);
     when "011011101000" => data <= triangle_rom(1768);
     when "011011101001" => data <= triangle_rom(1769);
     when "011011101010" => data <= triangle_rom(1770);
     when "011011101011" => data <= triangle_rom(1771);
     when "011011101100" => data <= triangle_rom(1772);
     when "011011101101" => data <= triangle_rom(1773);
     when "011011101110" => data <= triangle_rom(1774);
     when "011011101111" => data <= triangle_rom(1775);
     when "011011110000" => data <= triangle_rom(1776);
     when "011011110001" => data <= triangle_rom(1777);
     when "011011110010" => data <= triangle_rom(1778);
     when "011011110011" => data <= triangle_rom(1779);
     when "011011110100" => data <= triangle_rom(1780);
     when "011011110101" => data <= triangle_rom(1781);
     when "011011110110" => data <= triangle_rom(1782);
     when "011011110111" => data <= triangle_rom(1783);
     when "011011111000" => data <= triangle_rom(1784);
     when "011011111001" => data <= triangle_rom(1785);
     when "011011111010" => data <= triangle_rom(1786);
     when "011011111011" => data <= triangle_rom(1787);
     when "011011111100" => data <= triangle_rom(1788);
     when "011011111101" => data <= triangle_rom(1789);
     when "011011111110" => data <= triangle_rom(1790);
     when "011011111111" => data <= triangle_rom(1791);
     when "011100000000" => data <= triangle_rom(1792);
     when "011100000001" => data <= triangle_rom(1793);
     when "011100000010" => data <= triangle_rom(1794);
     when "011100000011" => data <= triangle_rom(1795);
     when "011100000100" => data <= triangle_rom(1796);
     when "011100000101" => data <= triangle_rom(1797);
     when "011100000110" => data <= triangle_rom(1798);
     when "011100000111" => data <= triangle_rom(1799);
     when "011100001000" => data <= triangle_rom(1800);
     when "011100001001" => data <= triangle_rom(1801);
     when "011100001010" => data <= triangle_rom(1802);
     when "011100001011" => data <= triangle_rom(1803);
     when "011100001100" => data <= triangle_rom(1804);
     when "011100001101" => data <= triangle_rom(1805);
     when "011100001110" => data <= triangle_rom(1806);
     when "011100001111" => data <= triangle_rom(1807);
     when "011100010000" => data <= triangle_rom(1808);
     when "011100010001" => data <= triangle_rom(1809);
     when "011100010010" => data <= triangle_rom(1810);
     when "011100010011" => data <= triangle_rom(1811);
     when "011100010100" => data <= triangle_rom(1812);
     when "011100010101" => data <= triangle_rom(1813);
     when "011100010110" => data <= triangle_rom(1814);
     when "011100010111" => data <= triangle_rom(1815);
     when "011100011000" => data <= triangle_rom(1816);
     when "011100011001" => data <= triangle_rom(1817);
     when "011100011010" => data <= triangle_rom(1818);
     when "011100011011" => data <= triangle_rom(1819);
     when "011100011100" => data <= triangle_rom(1820);
     when "011100011101" => data <= triangle_rom(1821);
     when "011100011110" => data <= triangle_rom(1822);
     when "011100011111" => data <= triangle_rom(1823);
     when "011100100000" => data <= triangle_rom(1824);
     when "011100100001" => data <= triangle_rom(1825);
     when "011100100010" => data <= triangle_rom(1826);
     when "011100100011" => data <= triangle_rom(1827);
     when "011100100100" => data <= triangle_rom(1828);
     when "011100100101" => data <= triangle_rom(1829);
     when "011100100110" => data <= triangle_rom(1830);
     when "011100100111" => data <= triangle_rom(1831);
     when "011100101000" => data <= triangle_rom(1832);
     when "011100101001" => data <= triangle_rom(1833);
     when "011100101010" => data <= triangle_rom(1834);
     when "011100101011" => data <= triangle_rom(1835);
     when "011100101100" => data <= triangle_rom(1836);
     when "011100101101" => data <= triangle_rom(1837);
     when "011100101110" => data <= triangle_rom(1838);
     when "011100101111" => data <= triangle_rom(1839);
     when "011100110000" => data <= triangle_rom(1840);
     when "011100110001" => data <= triangle_rom(1841);
     when "011100110010" => data <= triangle_rom(1842);
     when "011100110011" => data <= triangle_rom(1843);
     when "011100110100" => data <= triangle_rom(1844);
     when "011100110101" => data <= triangle_rom(1845);
     when "011100110110" => data <= triangle_rom(1846);
     when "011100110111" => data <= triangle_rom(1847);
     when "011100111000" => data <= triangle_rom(1848);
     when "011100111001" => data <= triangle_rom(1849);
     when "011100111010" => data <= triangle_rom(1850);
     when "011100111011" => data <= triangle_rom(1851);
     when "011100111100" => data <= triangle_rom(1852);
     when "011100111101" => data <= triangle_rom(1853);
     when "011100111110" => data <= triangle_rom(1854);
     when "011100111111" => data <= triangle_rom(1855);
     when "011101000000" => data <= triangle_rom(1856);
     when "011101000001" => data <= triangle_rom(1857);
     when "011101000010" => data <= triangle_rom(1858);
     when "011101000011" => data <= triangle_rom(1859);
     when "011101000100" => data <= triangle_rom(1860);
     when "011101000101" => data <= triangle_rom(1861);
     when "011101000110" => data <= triangle_rom(1862);
     when "011101000111" => data <= triangle_rom(1863);
     when "011101001000" => data <= triangle_rom(1864);
     when "011101001001" => data <= triangle_rom(1865);
     when "011101001010" => data <= triangle_rom(1866);
     when "011101001011" => data <= triangle_rom(1867);
     when "011101001100" => data <= triangle_rom(1868);
     when "011101001101" => data <= triangle_rom(1869);
     when "011101001110" => data <= triangle_rom(1870);
     when "011101001111" => data <= triangle_rom(1871);
     when "011101010000" => data <= triangle_rom(1872);
     when "011101010001" => data <= triangle_rom(1873);
     when "011101010010" => data <= triangle_rom(1874);
     when "011101010011" => data <= triangle_rom(1875);
     when "011101010100" => data <= triangle_rom(1876);
     when "011101010101" => data <= triangle_rom(1877);
     when "011101010110" => data <= triangle_rom(1878);
     when "011101010111" => data <= triangle_rom(1879);
     when "011101011000" => data <= triangle_rom(1880);
     when "011101011001" => data <= triangle_rom(1881);
     when "011101011010" => data <= triangle_rom(1882);
     when "011101011011" => data <= triangle_rom(1883);
     when "011101011100" => data <= triangle_rom(1884);
     when "011101011101" => data <= triangle_rom(1885);
     when "011101011110" => data <= triangle_rom(1886);
     when "011101011111" => data <= triangle_rom(1887);
     when "011101100000" => data <= triangle_rom(1888);
     when "011101100001" => data <= triangle_rom(1889);
     when "011101100010" => data <= triangle_rom(1890);
     when "011101100011" => data <= triangle_rom(1891);
     when "011101100100" => data <= triangle_rom(1892);
     when "011101100101" => data <= triangle_rom(1893);
     when "011101100110" => data <= triangle_rom(1894);
     when "011101100111" => data <= triangle_rom(1895);
     when "011101101000" => data <= triangle_rom(1896);
     when "011101101001" => data <= triangle_rom(1897);
     when "011101101010" => data <= triangle_rom(1898);
     when "011101101011" => data <= triangle_rom(1899);
     when "011101101100" => data <= triangle_rom(1900);
     when "011101101101" => data <= triangle_rom(1901);
     when "011101101110" => data <= triangle_rom(1902);
     when "011101101111" => data <= triangle_rom(1903);
     when "011101110000" => data <= triangle_rom(1904);
     when "011101110001" => data <= triangle_rom(1905);
     when "011101110010" => data <= triangle_rom(1906);
     when "011101110011" => data <= triangle_rom(1907);
     when "011101110100" => data <= triangle_rom(1908);
     when "011101110101" => data <= triangle_rom(1909);
     when "011101110110" => data <= triangle_rom(1910);
     when "011101110111" => data <= triangle_rom(1911);
     when "011101111000" => data <= triangle_rom(1912);
     when "011101111001" => data <= triangle_rom(1913);
     when "011101111010" => data <= triangle_rom(1914);
     when "011101111011" => data <= triangle_rom(1915);
     when "011101111100" => data <= triangle_rom(1916);
     when "011101111101" => data <= triangle_rom(1917);
     when "011101111110" => data <= triangle_rom(1918);
     when "011101111111" => data <= triangle_rom(1919);
     when "011110000000" => data <= triangle_rom(1920);
     when "011110000001" => data <= triangle_rom(1921);
     when "011110000010" => data <= triangle_rom(1922);
     when "011110000011" => data <= triangle_rom(1923);
     when "011110000100" => data <= triangle_rom(1924);
     when "011110000101" => data <= triangle_rom(1925);
     when "011110000110" => data <= triangle_rom(1926);
     when "011110000111" => data <= triangle_rom(1927);
     when "011110001000" => data <= triangle_rom(1928);
     when "011110001001" => data <= triangle_rom(1929);
     when "011110001010" => data <= triangle_rom(1930);
     when "011110001011" => data <= triangle_rom(1931);
     when "011110001100" => data <= triangle_rom(1932);
     when "011110001101" => data <= triangle_rom(1933);
     when "011110001110" => data <= triangle_rom(1934);
     when "011110001111" => data <= triangle_rom(1935);
     when "011110010000" => data <= triangle_rom(1936);
     when "011110010001" => data <= triangle_rom(1937);
     when "011110010010" => data <= triangle_rom(1938);
     when "011110010011" => data <= triangle_rom(1939);
     when "011110010100" => data <= triangle_rom(1940);
     when "011110010101" => data <= triangle_rom(1941);
     when "011110010110" => data <= triangle_rom(1942);
     when "011110010111" => data <= triangle_rom(1943);
     when "011110011000" => data <= triangle_rom(1944);
     when "011110011001" => data <= triangle_rom(1945);
     when "011110011010" => data <= triangle_rom(1946);
     when "011110011011" => data <= triangle_rom(1947);
     when "011110011100" => data <= triangle_rom(1948);
     when "011110011101" => data <= triangle_rom(1949);
     when "011110011110" => data <= triangle_rom(1950);
     when "011110011111" => data <= triangle_rom(1951);
     when "011110100000" => data <= triangle_rom(1952);
     when "011110100001" => data <= triangle_rom(1953);
     when "011110100010" => data <= triangle_rom(1954);
     when "011110100011" => data <= triangle_rom(1955);
     when "011110100100" => data <= triangle_rom(1956);
     when "011110100101" => data <= triangle_rom(1957);
     when "011110100110" => data <= triangle_rom(1958);
     when "011110100111" => data <= triangle_rom(1959);
     when "011110101000" => data <= triangle_rom(1960);
     when "011110101001" => data <= triangle_rom(1961);
     when "011110101010" => data <= triangle_rom(1962);
     when "011110101011" => data <= triangle_rom(1963);
     when "011110101100" => data <= triangle_rom(1964);
     when "011110101101" => data <= triangle_rom(1965);
     when "011110101110" => data <= triangle_rom(1966);
     when "011110101111" => data <= triangle_rom(1967);
     when "011110110000" => data <= triangle_rom(1968);
     when "011110110001" => data <= triangle_rom(1969);
     when "011110110010" => data <= triangle_rom(1970);
     when "011110110011" => data <= triangle_rom(1971);
     when "011110110100" => data <= triangle_rom(1972);
     when "011110110101" => data <= triangle_rom(1973);
     when "011110110110" => data <= triangle_rom(1974);
     when "011110110111" => data <= triangle_rom(1975);
     when "011110111000" => data <= triangle_rom(1976);
     when "011110111001" => data <= triangle_rom(1977);
     when "011110111010" => data <= triangle_rom(1978);
     when "011110111011" => data <= triangle_rom(1979);
     when "011110111100" => data <= triangle_rom(1980);
     when "011110111101" => data <= triangle_rom(1981);
     when "011110111110" => data <= triangle_rom(1982);
     when "011110111111" => data <= triangle_rom(1983);
     when "011111000000" => data <= triangle_rom(1984);
     when "011111000001" => data <= triangle_rom(1985);
     when "011111000010" => data <= triangle_rom(1986);
     when "011111000011" => data <= triangle_rom(1987);
     when "011111000100" => data <= triangle_rom(1988);
     when "011111000101" => data <= triangle_rom(1989);
     when "011111000110" => data <= triangle_rom(1990);
     when "011111000111" => data <= triangle_rom(1991);
     when "011111001000" => data <= triangle_rom(1992);
     when "011111001001" => data <= triangle_rom(1993);
     when "011111001010" => data <= triangle_rom(1994);
     when "011111001011" => data <= triangle_rom(1995);
     when "011111001100" => data <= triangle_rom(1996);
     when "011111001101" => data <= triangle_rom(1997);
     when "011111001110" => data <= triangle_rom(1998);
     when "011111001111" => data <= triangle_rom(1999);
     when "011111010000" => data <= triangle_rom(2000);
     when "011111010001" => data <= triangle_rom(2001);
     when "011111010010" => data <= triangle_rom(2002);
     when "011111010011" => data <= triangle_rom(2003);
     when "011111010100" => data <= triangle_rom(2004);
     when "011111010101" => data <= triangle_rom(2005);
     when "011111010110" => data <= triangle_rom(2006);
     when "011111010111" => data <= triangle_rom(2007);
     when "011111011000" => data <= triangle_rom(2008);
     when "011111011001" => data <= triangle_rom(2009);
     when "011111011010" => data <= triangle_rom(2010);
     when "011111011011" => data <= triangle_rom(2011);
     when "011111011100" => data <= triangle_rom(2012);
     when "011111011101" => data <= triangle_rom(2013);
     when "011111011110" => data <= triangle_rom(2014);
     when "011111011111" => data <= triangle_rom(2015);
     when "011111100000" => data <= triangle_rom(2016);
     when "011111100001" => data <= triangle_rom(2017);
     when "011111100010" => data <= triangle_rom(2018);
     when "011111100011" => data <= triangle_rom(2019);
     when "011111100100" => data <= triangle_rom(2020);
     when "011111100101" => data <= triangle_rom(2021);
     when "011111100110" => data <= triangle_rom(2022);
     when "011111100111" => data <= triangle_rom(2023);
     when "011111101000" => data <= triangle_rom(2024);
     when "011111101001" => data <= triangle_rom(2025);
     when "011111101010" => data <= triangle_rom(2026);
     when "011111101011" => data <= triangle_rom(2027);
     when "011111101100" => data <= triangle_rom(2028);
     when "011111101101" => data <= triangle_rom(2029);
     when "011111101110" => data <= triangle_rom(2030);
     when "011111101111" => data <= triangle_rom(2031);
     when "011111110000" => data <= triangle_rom(2032);
     when "011111110001" => data <= triangle_rom(2033);
     when "011111110010" => data <= triangle_rom(2034);
     when "011111110011" => data <= triangle_rom(2035);
     when "011111110100" => data <= triangle_rom(2036);
     when "011111110101" => data <= triangle_rom(2037);
     when "011111110110" => data <= triangle_rom(2038);
     when "011111110111" => data <= triangle_rom(2039);
     when "011111111000" => data <= triangle_rom(2040);
     when "011111111001" => data <= triangle_rom(2041);
     when "011111111010" => data <= triangle_rom(2042);
     when "011111111011" => data <= triangle_rom(2043);
     when "011111111100" => data <= triangle_rom(2044);
     when "011111111101" => data <= triangle_rom(2045);
     when "011111111110" => data <= triangle_rom(2046);
     when "011111111111" => data <= triangle_rom(2047);
     when "100000000000" => data <= triangle_rom(2048);
     when "100000000001" => data <= triangle_rom(2049);
     when "100000000010" => data <= triangle_rom(2050);
     when "100000000011" => data <= triangle_rom(2051);
     when "100000000100" => data <= triangle_rom(2052);
     when "100000000101" => data <= triangle_rom(2053);
     when "100000000110" => data <= triangle_rom(2054);
     when "100000000111" => data <= triangle_rom(2055);
     when "100000001000" => data <= triangle_rom(2056);
     when "100000001001" => data <= triangle_rom(2057);
     when "100000001010" => data <= triangle_rom(2058);
     when "100000001011" => data <= triangle_rom(2059);
     when "100000001100" => data <= triangle_rom(2060);
     when "100000001101" => data <= triangle_rom(2061);
     when "100000001110" => data <= triangle_rom(2062);
     when "100000001111" => data <= triangle_rom(2063);
     when "100000010000" => data <= triangle_rom(2064);
     when "100000010001" => data <= triangle_rom(2065);
     when "100000010010" => data <= triangle_rom(2066);
     when "100000010011" => data <= triangle_rom(2067);
     when "100000010100" => data <= triangle_rom(2068);
     when "100000010101" => data <= triangle_rom(2069);
     when "100000010110" => data <= triangle_rom(2070);
     when "100000010111" => data <= triangle_rom(2071);
     when "100000011000" => data <= triangle_rom(2072);
     when "100000011001" => data <= triangle_rom(2073);
     when "100000011010" => data <= triangle_rom(2074);
     when "100000011011" => data <= triangle_rom(2075);
     when "100000011100" => data <= triangle_rom(2076);
     when "100000011101" => data <= triangle_rom(2077);
     when "100000011110" => data <= triangle_rom(2078);
     when "100000011111" => data <= triangle_rom(2079);
     when "100000100000" => data <= triangle_rom(2080);
     when "100000100001" => data <= triangle_rom(2081);
     when "100000100010" => data <= triangle_rom(2082);
     when "100000100011" => data <= triangle_rom(2083);
     when "100000100100" => data <= triangle_rom(2084);
     when "100000100101" => data <= triangle_rom(2085);
     when "100000100110" => data <= triangle_rom(2086);
     when "100000100111" => data <= triangle_rom(2087);
     when "100000101000" => data <= triangle_rom(2088);
     when "100000101001" => data <= triangle_rom(2089);
     when "100000101010" => data <= triangle_rom(2090);
     when "100000101011" => data <= triangle_rom(2091);
     when "100000101100" => data <= triangle_rom(2092);
     when "100000101101" => data <= triangle_rom(2093);
     when "100000101110" => data <= triangle_rom(2094);
     when "100000101111" => data <= triangle_rom(2095);
     when "100000110000" => data <= triangle_rom(2096);
     when "100000110001" => data <= triangle_rom(2097);
     when "100000110010" => data <= triangle_rom(2098);
     when "100000110011" => data <= triangle_rom(2099);
     when "100000110100" => data <= triangle_rom(2100);
     when "100000110101" => data <= triangle_rom(2101);
     when "100000110110" => data <= triangle_rom(2102);
     when "100000110111" => data <= triangle_rom(2103);
     when "100000111000" => data <= triangle_rom(2104);
     when "100000111001" => data <= triangle_rom(2105);
     when "100000111010" => data <= triangle_rom(2106);
     when "100000111011" => data <= triangle_rom(2107);
     when "100000111100" => data <= triangle_rom(2108);
     when "100000111101" => data <= triangle_rom(2109);
     when "100000111110" => data <= triangle_rom(2110);
     when "100000111111" => data <= triangle_rom(2111);
     when "100001000000" => data <= triangle_rom(2112);
     when "100001000001" => data <= triangle_rom(2113);
     when "100001000010" => data <= triangle_rom(2114);
     when "100001000011" => data <= triangle_rom(2115);
     when "100001000100" => data <= triangle_rom(2116);
     when "100001000101" => data <= triangle_rom(2117);
     when "100001000110" => data <= triangle_rom(2118);
     when "100001000111" => data <= triangle_rom(2119);
     when "100001001000" => data <= triangle_rom(2120);
     when "100001001001" => data <= triangle_rom(2121);
     when "100001001010" => data <= triangle_rom(2122);
     when "100001001011" => data <= triangle_rom(2123);
     when "100001001100" => data <= triangle_rom(2124);
     when "100001001101" => data <= triangle_rom(2125);
     when "100001001110" => data <= triangle_rom(2126);
     when "100001001111" => data <= triangle_rom(2127);
     when "100001010000" => data <= triangle_rom(2128);
     when "100001010001" => data <= triangle_rom(2129);
     when "100001010010" => data <= triangle_rom(2130);
     when "100001010011" => data <= triangle_rom(2131);
     when "100001010100" => data <= triangle_rom(2132);
     when "100001010101" => data <= triangle_rom(2133);
     when "100001010110" => data <= triangle_rom(2134);
     when "100001010111" => data <= triangle_rom(2135);
     when "100001011000" => data <= triangle_rom(2136);
     when "100001011001" => data <= triangle_rom(2137);
     when "100001011010" => data <= triangle_rom(2138);
     when "100001011011" => data <= triangle_rom(2139);
     when "100001011100" => data <= triangle_rom(2140);
     when "100001011101" => data <= triangle_rom(2141);
     when "100001011110" => data <= triangle_rom(2142);
     when "100001011111" => data <= triangle_rom(2143);
     when "100001100000" => data <= triangle_rom(2144);
     when "100001100001" => data <= triangle_rom(2145);
     when "100001100010" => data <= triangle_rom(2146);
     when "100001100011" => data <= triangle_rom(2147);
     when "100001100100" => data <= triangle_rom(2148);
     when "100001100101" => data <= triangle_rom(2149);
     when "100001100110" => data <= triangle_rom(2150);
     when "100001100111" => data <= triangle_rom(2151);
     when "100001101000" => data <= triangle_rom(2152);
     when "100001101001" => data <= triangle_rom(2153);
     when "100001101010" => data <= triangle_rom(2154);
     when "100001101011" => data <= triangle_rom(2155);
     when "100001101100" => data <= triangle_rom(2156);
     when "100001101101" => data <= triangle_rom(2157);
     when "100001101110" => data <= triangle_rom(2158);
     when "100001101111" => data <= triangle_rom(2159);
     when "100001110000" => data <= triangle_rom(2160);
     when "100001110001" => data <= triangle_rom(2161);
     when "100001110010" => data <= triangle_rom(2162);
     when "100001110011" => data <= triangle_rom(2163);
     when "100001110100" => data <= triangle_rom(2164);
     when "100001110101" => data <= triangle_rom(2165);
     when "100001110110" => data <= triangle_rom(2166);
     when "100001110111" => data <= triangle_rom(2167);
     when "100001111000" => data <= triangle_rom(2168);
     when "100001111001" => data <= triangle_rom(2169);
     when "100001111010" => data <= triangle_rom(2170);
     when "100001111011" => data <= triangle_rom(2171);
     when "100001111100" => data <= triangle_rom(2172);
     when "100001111101" => data <= triangle_rom(2173);
     when "100001111110" => data <= triangle_rom(2174);
     when "100001111111" => data <= triangle_rom(2175);
     when "100010000000" => data <= triangle_rom(2176);
     when "100010000001" => data <= triangle_rom(2177);
     when "100010000010" => data <= triangle_rom(2178);
     when "100010000011" => data <= triangle_rom(2179);
     when "100010000100" => data <= triangle_rom(2180);
     when "100010000101" => data <= triangle_rom(2181);
     when "100010000110" => data <= triangle_rom(2182);
     when "100010000111" => data <= triangle_rom(2183);
     when "100010001000" => data <= triangle_rom(2184);
     when "100010001001" => data <= triangle_rom(2185);
     when "100010001010" => data <= triangle_rom(2186);
     when "100010001011" => data <= triangle_rom(2187);
     when "100010001100" => data <= triangle_rom(2188);
     when "100010001101" => data <= triangle_rom(2189);
     when "100010001110" => data <= triangle_rom(2190);
     when "100010001111" => data <= triangle_rom(2191);
     when "100010010000" => data <= triangle_rom(2192);
     when "100010010001" => data <= triangle_rom(2193);
     when "100010010010" => data <= triangle_rom(2194);
     when "100010010011" => data <= triangle_rom(2195);
     when "100010010100" => data <= triangle_rom(2196);
     when "100010010101" => data <= triangle_rom(2197);
     when "100010010110" => data <= triangle_rom(2198);
     when "100010010111" => data <= triangle_rom(2199);
     when "100010011000" => data <= triangle_rom(2200);
     when "100010011001" => data <= triangle_rom(2201);
     when "100010011010" => data <= triangle_rom(2202);
     when "100010011011" => data <= triangle_rom(2203);
     when "100010011100" => data <= triangle_rom(2204);
     when "100010011101" => data <= triangle_rom(2205);
     when "100010011110" => data <= triangle_rom(2206);
     when "100010011111" => data <= triangle_rom(2207);
     when "100010100000" => data <= triangle_rom(2208);
     when "100010100001" => data <= triangle_rom(2209);
     when "100010100010" => data <= triangle_rom(2210);
     when "100010100011" => data <= triangle_rom(2211);
     when "100010100100" => data <= triangle_rom(2212);
     when "100010100101" => data <= triangle_rom(2213);
     when "100010100110" => data <= triangle_rom(2214);
     when "100010100111" => data <= triangle_rom(2215);
     when "100010101000" => data <= triangle_rom(2216);
     when "100010101001" => data <= triangle_rom(2217);
     when "100010101010" => data <= triangle_rom(2218);
     when "100010101011" => data <= triangle_rom(2219);
     when "100010101100" => data <= triangle_rom(2220);
     when "100010101101" => data <= triangle_rom(2221);
     when "100010101110" => data <= triangle_rom(2222);
     when "100010101111" => data <= triangle_rom(2223);
     when "100010110000" => data <= triangle_rom(2224);
     when "100010110001" => data <= triangle_rom(2225);
     when "100010110010" => data <= triangle_rom(2226);
     when "100010110011" => data <= triangle_rom(2227);
     when "100010110100" => data <= triangle_rom(2228);
     when "100010110101" => data <= triangle_rom(2229);
     when "100010110110" => data <= triangle_rom(2230);
     when "100010110111" => data <= triangle_rom(2231);
     when "100010111000" => data <= triangle_rom(2232);
     when "100010111001" => data <= triangle_rom(2233);
     when "100010111010" => data <= triangle_rom(2234);
     when "100010111011" => data <= triangle_rom(2235);
     when "100010111100" => data <= triangle_rom(2236);
     when "100010111101" => data <= triangle_rom(2237);
     when "100010111110" => data <= triangle_rom(2238);
     when "100010111111" => data <= triangle_rom(2239);
     when "100011000000" => data <= triangle_rom(2240);
     when "100011000001" => data <= triangle_rom(2241);
     when "100011000010" => data <= triangle_rom(2242);
     when "100011000011" => data <= triangle_rom(2243);
     when "100011000100" => data <= triangle_rom(2244);
     when "100011000101" => data <= triangle_rom(2245);
     when "100011000110" => data <= triangle_rom(2246);
     when "100011000111" => data <= triangle_rom(2247);
     when "100011001000" => data <= triangle_rom(2248);
     when "100011001001" => data <= triangle_rom(2249);
     when "100011001010" => data <= triangle_rom(2250);
     when "100011001011" => data <= triangle_rom(2251);
     when "100011001100" => data <= triangle_rom(2252);
     when "100011001101" => data <= triangle_rom(2253);
     when "100011001110" => data <= triangle_rom(2254);
     when "100011001111" => data <= triangle_rom(2255);
     when "100011010000" => data <= triangle_rom(2256);
     when "100011010001" => data <= triangle_rom(2257);
     when "100011010010" => data <= triangle_rom(2258);
     when "100011010011" => data <= triangle_rom(2259);
     when "100011010100" => data <= triangle_rom(2260);
     when "100011010101" => data <= triangle_rom(2261);
     when "100011010110" => data <= triangle_rom(2262);
     when "100011010111" => data <= triangle_rom(2263);
     when "100011011000" => data <= triangle_rom(2264);
     when "100011011001" => data <= triangle_rom(2265);
     when "100011011010" => data <= triangle_rom(2266);
     when "100011011011" => data <= triangle_rom(2267);
     when "100011011100" => data <= triangle_rom(2268);
     when "100011011101" => data <= triangle_rom(2269);
     when "100011011110" => data <= triangle_rom(2270);
     when "100011011111" => data <= triangle_rom(2271);
     when "100011100000" => data <= triangle_rom(2272);
     when "100011100001" => data <= triangle_rom(2273);
     when "100011100010" => data <= triangle_rom(2274);
     when "100011100011" => data <= triangle_rom(2275);
     when "100011100100" => data <= triangle_rom(2276);
     when "100011100101" => data <= triangle_rom(2277);
     when "100011100110" => data <= triangle_rom(2278);
     when "100011100111" => data <= triangle_rom(2279);
     when "100011101000" => data <= triangle_rom(2280);
     when "100011101001" => data <= triangle_rom(2281);
     when "100011101010" => data <= triangle_rom(2282);
     when "100011101011" => data <= triangle_rom(2283);
     when "100011101100" => data <= triangle_rom(2284);
     when "100011101101" => data <= triangle_rom(2285);
     when "100011101110" => data <= triangle_rom(2286);
     when "100011101111" => data <= triangle_rom(2287);
     when "100011110000" => data <= triangle_rom(2288);
     when "100011110001" => data <= triangle_rom(2289);
     when "100011110010" => data <= triangle_rom(2290);
     when "100011110011" => data <= triangle_rom(2291);
     when "100011110100" => data <= triangle_rom(2292);
     when "100011110101" => data <= triangle_rom(2293);
     when "100011110110" => data <= triangle_rom(2294);
     when "100011110111" => data <= triangle_rom(2295);
     when "100011111000" => data <= triangle_rom(2296);
     when "100011111001" => data <= triangle_rom(2297);
     when "100011111010" => data <= triangle_rom(2298);
     when "100011111011" => data <= triangle_rom(2299);
     when "100011111100" => data <= triangle_rom(2300);
     when "100011111101" => data <= triangle_rom(2301);
     when "100011111110" => data <= triangle_rom(2302);
     when "100011111111" => data <= triangle_rom(2303);
     when "100100000000" => data <= triangle_rom(2304);
     when "100100000001" => data <= triangle_rom(2305);
     when "100100000010" => data <= triangle_rom(2306);
     when "100100000011" => data <= triangle_rom(2307);
     when "100100000100" => data <= triangle_rom(2308);
     when "100100000101" => data <= triangle_rom(2309);
     when "100100000110" => data <= triangle_rom(2310);
     when "100100000111" => data <= triangle_rom(2311);
     when "100100001000" => data <= triangle_rom(2312);
     when "100100001001" => data <= triangle_rom(2313);
     when "100100001010" => data <= triangle_rom(2314);
     when "100100001011" => data <= triangle_rom(2315);
     when "100100001100" => data <= triangle_rom(2316);
     when "100100001101" => data <= triangle_rom(2317);
     when "100100001110" => data <= triangle_rom(2318);
     when "100100001111" => data <= triangle_rom(2319);
     when "100100010000" => data <= triangle_rom(2320);
     when "100100010001" => data <= triangle_rom(2321);
     when "100100010010" => data <= triangle_rom(2322);
     when "100100010011" => data <= triangle_rom(2323);
     when "100100010100" => data <= triangle_rom(2324);
     when "100100010101" => data <= triangle_rom(2325);
     when "100100010110" => data <= triangle_rom(2326);
     when "100100010111" => data <= triangle_rom(2327);
     when "100100011000" => data <= triangle_rom(2328);
     when "100100011001" => data <= triangle_rom(2329);
     when "100100011010" => data <= triangle_rom(2330);
     when "100100011011" => data <= triangle_rom(2331);
     when "100100011100" => data <= triangle_rom(2332);
     when "100100011101" => data <= triangle_rom(2333);
     when "100100011110" => data <= triangle_rom(2334);
     when "100100011111" => data <= triangle_rom(2335);
     when "100100100000" => data <= triangle_rom(2336);
     when "100100100001" => data <= triangle_rom(2337);
     when "100100100010" => data <= triangle_rom(2338);
     when "100100100011" => data <= triangle_rom(2339);
     when "100100100100" => data <= triangle_rom(2340);
     when "100100100101" => data <= triangle_rom(2341);
     when "100100100110" => data <= triangle_rom(2342);
     when "100100100111" => data <= triangle_rom(2343);
     when "100100101000" => data <= triangle_rom(2344);
     when "100100101001" => data <= triangle_rom(2345);
     when "100100101010" => data <= triangle_rom(2346);
     when "100100101011" => data <= triangle_rom(2347);
     when "100100101100" => data <= triangle_rom(2348);
     when "100100101101" => data <= triangle_rom(2349);
     when "100100101110" => data <= triangle_rom(2350);
     when "100100101111" => data <= triangle_rom(2351);
     when "100100110000" => data <= triangle_rom(2352);
     when "100100110001" => data <= triangle_rom(2353);
     when "100100110010" => data <= triangle_rom(2354);
     when "100100110011" => data <= triangle_rom(2355);
     when "100100110100" => data <= triangle_rom(2356);
     when "100100110101" => data <= triangle_rom(2357);
     when "100100110110" => data <= triangle_rom(2358);
     when "100100110111" => data <= triangle_rom(2359);
     when "100100111000" => data <= triangle_rom(2360);
     when "100100111001" => data <= triangle_rom(2361);
     when "100100111010" => data <= triangle_rom(2362);
     when "100100111011" => data <= triangle_rom(2363);
     when "100100111100" => data <= triangle_rom(2364);
     when "100100111101" => data <= triangle_rom(2365);
     when "100100111110" => data <= triangle_rom(2366);
     when "100100111111" => data <= triangle_rom(2367);
     when "100101000000" => data <= triangle_rom(2368);
     when "100101000001" => data <= triangle_rom(2369);
     when "100101000010" => data <= triangle_rom(2370);
     when "100101000011" => data <= triangle_rom(2371);
     when "100101000100" => data <= triangle_rom(2372);
     when "100101000101" => data <= triangle_rom(2373);
     when "100101000110" => data <= triangle_rom(2374);
     when "100101000111" => data <= triangle_rom(2375);
     when "100101001000" => data <= triangle_rom(2376);
     when "100101001001" => data <= triangle_rom(2377);
     when "100101001010" => data <= triangle_rom(2378);
     when "100101001011" => data <= triangle_rom(2379);
     when "100101001100" => data <= triangle_rom(2380);
     when "100101001101" => data <= triangle_rom(2381);
     when "100101001110" => data <= triangle_rom(2382);
     when "100101001111" => data <= triangle_rom(2383);
     when "100101010000" => data <= triangle_rom(2384);
     when "100101010001" => data <= triangle_rom(2385);
     when "100101010010" => data <= triangle_rom(2386);
     when "100101010011" => data <= triangle_rom(2387);
     when "100101010100" => data <= triangle_rom(2388);
     when "100101010101" => data <= triangle_rom(2389);
     when "100101010110" => data <= triangle_rom(2390);
     when "100101010111" => data <= triangle_rom(2391);
     when "100101011000" => data <= triangle_rom(2392);
     when "100101011001" => data <= triangle_rom(2393);
     when "100101011010" => data <= triangle_rom(2394);
     when "100101011011" => data <= triangle_rom(2395);
     when "100101011100" => data <= triangle_rom(2396);
     when "100101011101" => data <= triangle_rom(2397);
     when "100101011110" => data <= triangle_rom(2398);
     when "100101011111" => data <= triangle_rom(2399);
     when "100101100000" => data <= triangle_rom(2400);
     when "100101100001" => data <= triangle_rom(2401);
     when "100101100010" => data <= triangle_rom(2402);
     when "100101100011" => data <= triangle_rom(2403);
     when "100101100100" => data <= triangle_rom(2404);
     when "100101100101" => data <= triangle_rom(2405);
     when "100101100110" => data <= triangle_rom(2406);
     when "100101100111" => data <= triangle_rom(2407);
     when "100101101000" => data <= triangle_rom(2408);
     when "100101101001" => data <= triangle_rom(2409);
     when "100101101010" => data <= triangle_rom(2410);
     when "100101101011" => data <= triangle_rom(2411);
     when "100101101100" => data <= triangle_rom(2412);
     when "100101101101" => data <= triangle_rom(2413);
     when "100101101110" => data <= triangle_rom(2414);
     when "100101101111" => data <= triangle_rom(2415);
     when "100101110000" => data <= triangle_rom(2416);
     when "100101110001" => data <= triangle_rom(2417);
     when "100101110010" => data <= triangle_rom(2418);
     when "100101110011" => data <= triangle_rom(2419);
     when "100101110100" => data <= triangle_rom(2420);
     when "100101110101" => data <= triangle_rom(2421);
     when "100101110110" => data <= triangle_rom(2422);
     when "100101110111" => data <= triangle_rom(2423);
     when "100101111000" => data <= triangle_rom(2424);
     when "100101111001" => data <= triangle_rom(2425);
     when "100101111010" => data <= triangle_rom(2426);
     when "100101111011" => data <= triangle_rom(2427);
     when "100101111100" => data <= triangle_rom(2428);
     when "100101111101" => data <= triangle_rom(2429);
     when "100101111110" => data <= triangle_rom(2430);
     when "100101111111" => data <= triangle_rom(2431);
     when "100110000000" => data <= triangle_rom(2432);
     when "100110000001" => data <= triangle_rom(2433);
     when "100110000010" => data <= triangle_rom(2434);
     when "100110000011" => data <= triangle_rom(2435);
     when "100110000100" => data <= triangle_rom(2436);
     when "100110000101" => data <= triangle_rom(2437);
     when "100110000110" => data <= triangle_rom(2438);
     when "100110000111" => data <= triangle_rom(2439);
     when "100110001000" => data <= triangle_rom(2440);
     when "100110001001" => data <= triangle_rom(2441);
     when "100110001010" => data <= triangle_rom(2442);
     when "100110001011" => data <= triangle_rom(2443);
     when "100110001100" => data <= triangle_rom(2444);
     when "100110001101" => data <= triangle_rom(2445);
     when "100110001110" => data <= triangle_rom(2446);
     when "100110001111" => data <= triangle_rom(2447);
     when "100110010000" => data <= triangle_rom(2448);
     when "100110010001" => data <= triangle_rom(2449);
     when "100110010010" => data <= triangle_rom(2450);
     when "100110010011" => data <= triangle_rom(2451);
     when "100110010100" => data <= triangle_rom(2452);
     when "100110010101" => data <= triangle_rom(2453);
     when "100110010110" => data <= triangle_rom(2454);
     when "100110010111" => data <= triangle_rom(2455);
     when "100110011000" => data <= triangle_rom(2456);
     when "100110011001" => data <= triangle_rom(2457);
     when "100110011010" => data <= triangle_rom(2458);
     when "100110011011" => data <= triangle_rom(2459);
     when "100110011100" => data <= triangle_rom(2460);
     when "100110011101" => data <= triangle_rom(2461);
     when "100110011110" => data <= triangle_rom(2462);
     when "100110011111" => data <= triangle_rom(2463);
     when "100110100000" => data <= triangle_rom(2464);
     when "100110100001" => data <= triangle_rom(2465);
     when "100110100010" => data <= triangle_rom(2466);
     when "100110100011" => data <= triangle_rom(2467);
     when "100110100100" => data <= triangle_rom(2468);
     when "100110100101" => data <= triangle_rom(2469);
     when "100110100110" => data <= triangle_rom(2470);
     when "100110100111" => data <= triangle_rom(2471);
     when "100110101000" => data <= triangle_rom(2472);
     when "100110101001" => data <= triangle_rom(2473);
     when "100110101010" => data <= triangle_rom(2474);
     when "100110101011" => data <= triangle_rom(2475);
     when "100110101100" => data <= triangle_rom(2476);
     when "100110101101" => data <= triangle_rom(2477);
     when "100110101110" => data <= triangle_rom(2478);
     when "100110101111" => data <= triangle_rom(2479);
     when "100110110000" => data <= triangle_rom(2480);
     when "100110110001" => data <= triangle_rom(2481);
     when "100110110010" => data <= triangle_rom(2482);
     when "100110110011" => data <= triangle_rom(2483);
     when "100110110100" => data <= triangle_rom(2484);
     when "100110110101" => data <= triangle_rom(2485);
     when "100110110110" => data <= triangle_rom(2486);
     when "100110110111" => data <= triangle_rom(2487);
     when "100110111000" => data <= triangle_rom(2488);
     when "100110111001" => data <= triangle_rom(2489);
     when "100110111010" => data <= triangle_rom(2490);
     when "100110111011" => data <= triangle_rom(2491);
     when "100110111100" => data <= triangle_rom(2492);
     when "100110111101" => data <= triangle_rom(2493);
     when "100110111110" => data <= triangle_rom(2494);
     when "100110111111" => data <= triangle_rom(2495);
     when "100111000000" => data <= triangle_rom(2496);
     when "100111000001" => data <= triangle_rom(2497);
     when "100111000010" => data <= triangle_rom(2498);
     when "100111000011" => data <= triangle_rom(2499);
     when "100111000100" => data <= triangle_rom(2500);
     when "100111000101" => data <= triangle_rom(2501);
     when "100111000110" => data <= triangle_rom(2502);
     when "100111000111" => data <= triangle_rom(2503);
     when "100111001000" => data <= triangle_rom(2504);
     when "100111001001" => data <= triangle_rom(2505);
     when "100111001010" => data <= triangle_rom(2506);
     when "100111001011" => data <= triangle_rom(2507);
     when "100111001100" => data <= triangle_rom(2508);
     when "100111001101" => data <= triangle_rom(2509);
     when "100111001110" => data <= triangle_rom(2510);
     when "100111001111" => data <= triangle_rom(2511);
     when "100111010000" => data <= triangle_rom(2512);
     when "100111010001" => data <= triangle_rom(2513);
     when "100111010010" => data <= triangle_rom(2514);
     when "100111010011" => data <= triangle_rom(2515);
     when "100111010100" => data <= triangle_rom(2516);
     when "100111010101" => data <= triangle_rom(2517);
     when "100111010110" => data <= triangle_rom(2518);
     when "100111010111" => data <= triangle_rom(2519);
     when "100111011000" => data <= triangle_rom(2520);
     when "100111011001" => data <= triangle_rom(2521);
     when "100111011010" => data <= triangle_rom(2522);
     when "100111011011" => data <= triangle_rom(2523);
     when "100111011100" => data <= triangle_rom(2524);
     when "100111011101" => data <= triangle_rom(2525);
     when "100111011110" => data <= triangle_rom(2526);
     when "100111011111" => data <= triangle_rom(2527);
     when "100111100000" => data <= triangle_rom(2528);
     when "100111100001" => data <= triangle_rom(2529);
     when "100111100010" => data <= triangle_rom(2530);
     when "100111100011" => data <= triangle_rom(2531);
     when "100111100100" => data <= triangle_rom(2532);
     when "100111100101" => data <= triangle_rom(2533);
     when "100111100110" => data <= triangle_rom(2534);
     when "100111100111" => data <= triangle_rom(2535);
     when "100111101000" => data <= triangle_rom(2536);
     when "100111101001" => data <= triangle_rom(2537);
     when "100111101010" => data <= triangle_rom(2538);
     when "100111101011" => data <= triangle_rom(2539);
     when "100111101100" => data <= triangle_rom(2540);
     when "100111101101" => data <= triangle_rom(2541);
     when "100111101110" => data <= triangle_rom(2542);
     when "100111101111" => data <= triangle_rom(2543);
     when "100111110000" => data <= triangle_rom(2544);
     when "100111110001" => data <= triangle_rom(2545);
     when "100111110010" => data <= triangle_rom(2546);
     when "100111110011" => data <= triangle_rom(2547);
     when "100111110100" => data <= triangle_rom(2548);
     when "100111110101" => data <= triangle_rom(2549);
     when "100111110110" => data <= triangle_rom(2550);
     when "100111110111" => data <= triangle_rom(2551);
     when "100111111000" => data <= triangle_rom(2552);
     when "100111111001" => data <= triangle_rom(2553);
     when "100111111010" => data <= triangle_rom(2554);
     when "100111111011" => data <= triangle_rom(2555);
     when "100111111100" => data <= triangle_rom(2556);
     when "100111111101" => data <= triangle_rom(2557);
     when "100111111110" => data <= triangle_rom(2558);
     when "100111111111" => data <= triangle_rom(2559);
     when "101000000000" => data <= triangle_rom(2560);
     when "101000000001" => data <= triangle_rom(2561);
     when "101000000010" => data <= triangle_rom(2562);
     when "101000000011" => data <= triangle_rom(2563);
     when "101000000100" => data <= triangle_rom(2564);
     when "101000000101" => data <= triangle_rom(2565);
     when "101000000110" => data <= triangle_rom(2566);
     when "101000000111" => data <= triangle_rom(2567);
     when "101000001000" => data <= triangle_rom(2568);
     when "101000001001" => data <= triangle_rom(2569);
     when "101000001010" => data <= triangle_rom(2570);
     when "101000001011" => data <= triangle_rom(2571);
     when "101000001100" => data <= triangle_rom(2572);
     when "101000001101" => data <= triangle_rom(2573);
     when "101000001110" => data <= triangle_rom(2574);
     when "101000001111" => data <= triangle_rom(2575);
     when "101000010000" => data <= triangle_rom(2576);
     when "101000010001" => data <= triangle_rom(2577);
     when "101000010010" => data <= triangle_rom(2578);
     when "101000010011" => data <= triangle_rom(2579);
     when "101000010100" => data <= triangle_rom(2580);
     when "101000010101" => data <= triangle_rom(2581);
     when "101000010110" => data <= triangle_rom(2582);
     when "101000010111" => data <= triangle_rom(2583);
     when "101000011000" => data <= triangle_rom(2584);
     when "101000011001" => data <= triangle_rom(2585);
     when "101000011010" => data <= triangle_rom(2586);
     when "101000011011" => data <= triangle_rom(2587);
     when "101000011100" => data <= triangle_rom(2588);
     when "101000011101" => data <= triangle_rom(2589);
     when "101000011110" => data <= triangle_rom(2590);
     when "101000011111" => data <= triangle_rom(2591);
     when "101000100000" => data <= triangle_rom(2592);
     when "101000100001" => data <= triangle_rom(2593);
     when "101000100010" => data <= triangle_rom(2594);
     when "101000100011" => data <= triangle_rom(2595);
     when "101000100100" => data <= triangle_rom(2596);
     when "101000100101" => data <= triangle_rom(2597);
     when "101000100110" => data <= triangle_rom(2598);
     when "101000100111" => data <= triangle_rom(2599);
     when "101000101000" => data <= triangle_rom(2600);
     when "101000101001" => data <= triangle_rom(2601);
     when "101000101010" => data <= triangle_rom(2602);
     when "101000101011" => data <= triangle_rom(2603);
     when "101000101100" => data <= triangle_rom(2604);
     when "101000101101" => data <= triangle_rom(2605);
     when "101000101110" => data <= triangle_rom(2606);
     when "101000101111" => data <= triangle_rom(2607);
     when "101000110000" => data <= triangle_rom(2608);
     when "101000110001" => data <= triangle_rom(2609);
     when "101000110010" => data <= triangle_rom(2610);
     when "101000110011" => data <= triangle_rom(2611);
     when "101000110100" => data <= triangle_rom(2612);
     when "101000110101" => data <= triangle_rom(2613);
     when "101000110110" => data <= triangle_rom(2614);
     when "101000110111" => data <= triangle_rom(2615);
     when "101000111000" => data <= triangle_rom(2616);
     when "101000111001" => data <= triangle_rom(2617);
     when "101000111010" => data <= triangle_rom(2618);
     when "101000111011" => data <= triangle_rom(2619);
     when "101000111100" => data <= triangle_rom(2620);
     when "101000111101" => data <= triangle_rom(2621);
     when "101000111110" => data <= triangle_rom(2622);
     when "101000111111" => data <= triangle_rom(2623);
     when "101001000000" => data <= triangle_rom(2624);
     when "101001000001" => data <= triangle_rom(2625);
     when "101001000010" => data <= triangle_rom(2626);
     when "101001000011" => data <= triangle_rom(2627);
     when "101001000100" => data <= triangle_rom(2628);
     when "101001000101" => data <= triangle_rom(2629);
     when "101001000110" => data <= triangle_rom(2630);
     when "101001000111" => data <= triangle_rom(2631);
     when "101001001000" => data <= triangle_rom(2632);
     when "101001001001" => data <= triangle_rom(2633);
     when "101001001010" => data <= triangle_rom(2634);
     when "101001001011" => data <= triangle_rom(2635);
     when "101001001100" => data <= triangle_rom(2636);
     when "101001001101" => data <= triangle_rom(2637);
     when "101001001110" => data <= triangle_rom(2638);
     when "101001001111" => data <= triangle_rom(2639);
     when "101001010000" => data <= triangle_rom(2640);
     when "101001010001" => data <= triangle_rom(2641);
     when "101001010010" => data <= triangle_rom(2642);
     when "101001010011" => data <= triangle_rom(2643);
     when "101001010100" => data <= triangle_rom(2644);
     when "101001010101" => data <= triangle_rom(2645);
     when "101001010110" => data <= triangle_rom(2646);
     when "101001010111" => data <= triangle_rom(2647);
     when "101001011000" => data <= triangle_rom(2648);
     when "101001011001" => data <= triangle_rom(2649);
     when "101001011010" => data <= triangle_rom(2650);
     when "101001011011" => data <= triangle_rom(2651);
     when "101001011100" => data <= triangle_rom(2652);
     when "101001011101" => data <= triangle_rom(2653);
     when "101001011110" => data <= triangle_rom(2654);
     when "101001011111" => data <= triangle_rom(2655);
     when "101001100000" => data <= triangle_rom(2656);
     when "101001100001" => data <= triangle_rom(2657);
     when "101001100010" => data <= triangle_rom(2658);
     when "101001100011" => data <= triangle_rom(2659);
     when "101001100100" => data <= triangle_rom(2660);
     when "101001100101" => data <= triangle_rom(2661);
     when "101001100110" => data <= triangle_rom(2662);
     when "101001100111" => data <= triangle_rom(2663);
     when "101001101000" => data <= triangle_rom(2664);
     when "101001101001" => data <= triangle_rom(2665);
     when "101001101010" => data <= triangle_rom(2666);
     when "101001101011" => data <= triangle_rom(2667);
     when "101001101100" => data <= triangle_rom(2668);
     when "101001101101" => data <= triangle_rom(2669);
     when "101001101110" => data <= triangle_rom(2670);
     when "101001101111" => data <= triangle_rom(2671);
     when "101001110000" => data <= triangle_rom(2672);
     when "101001110001" => data <= triangle_rom(2673);
     when "101001110010" => data <= triangle_rom(2674);
     when "101001110011" => data <= triangle_rom(2675);
     when "101001110100" => data <= triangle_rom(2676);
     when "101001110101" => data <= triangle_rom(2677);
     when "101001110110" => data <= triangle_rom(2678);
     when "101001110111" => data <= triangle_rom(2679);
     when "101001111000" => data <= triangle_rom(2680);
     when "101001111001" => data <= triangle_rom(2681);
     when "101001111010" => data <= triangle_rom(2682);
     when "101001111011" => data <= triangle_rom(2683);
     when "101001111100" => data <= triangle_rom(2684);
     when "101001111101" => data <= triangle_rom(2685);
     when "101001111110" => data <= triangle_rom(2686);
     when "101001111111" => data <= triangle_rom(2687);
     when "101010000000" => data <= triangle_rom(2688);
     when "101010000001" => data <= triangle_rom(2689);
     when "101010000010" => data <= triangle_rom(2690);
     when "101010000011" => data <= triangle_rom(2691);
     when "101010000100" => data <= triangle_rom(2692);
     when "101010000101" => data <= triangle_rom(2693);
     when "101010000110" => data <= triangle_rom(2694);
     when "101010000111" => data <= triangle_rom(2695);
     when "101010001000" => data <= triangle_rom(2696);
     when "101010001001" => data <= triangle_rom(2697);
     when "101010001010" => data <= triangle_rom(2698);
     when "101010001011" => data <= triangle_rom(2699);
     when "101010001100" => data <= triangle_rom(2700);
     when "101010001101" => data <= triangle_rom(2701);
     when "101010001110" => data <= triangle_rom(2702);
     when "101010001111" => data <= triangle_rom(2703);
     when "101010010000" => data <= triangle_rom(2704);
     when "101010010001" => data <= triangle_rom(2705);
     when "101010010010" => data <= triangle_rom(2706);
     when "101010010011" => data <= triangle_rom(2707);
     when "101010010100" => data <= triangle_rom(2708);
     when "101010010101" => data <= triangle_rom(2709);
     when "101010010110" => data <= triangle_rom(2710);
     when "101010010111" => data <= triangle_rom(2711);
     when "101010011000" => data <= triangle_rom(2712);
     when "101010011001" => data <= triangle_rom(2713);
     when "101010011010" => data <= triangle_rom(2714);
     when "101010011011" => data <= triangle_rom(2715);
     when "101010011100" => data <= triangle_rom(2716);
     when "101010011101" => data <= triangle_rom(2717);
     when "101010011110" => data <= triangle_rom(2718);
     when "101010011111" => data <= triangle_rom(2719);
     when "101010100000" => data <= triangle_rom(2720);
     when "101010100001" => data <= triangle_rom(2721);
     when "101010100010" => data <= triangle_rom(2722);
     when "101010100011" => data <= triangle_rom(2723);
     when "101010100100" => data <= triangle_rom(2724);
     when "101010100101" => data <= triangle_rom(2725);
     when "101010100110" => data <= triangle_rom(2726);
     when "101010100111" => data <= triangle_rom(2727);
     when "101010101000" => data <= triangle_rom(2728);
     when "101010101001" => data <= triangle_rom(2729);
     when "101010101010" => data <= triangle_rom(2730);
     when "101010101011" => data <= triangle_rom(2731);
     when "101010101100" => data <= triangle_rom(2732);
     when "101010101101" => data <= triangle_rom(2733);
     when "101010101110" => data <= triangle_rom(2734);
     when "101010101111" => data <= triangle_rom(2735);
     when "101010110000" => data <= triangle_rom(2736);
     when "101010110001" => data <= triangle_rom(2737);
     when "101010110010" => data <= triangle_rom(2738);
     when "101010110011" => data <= triangle_rom(2739);
     when "101010110100" => data <= triangle_rom(2740);
     when "101010110101" => data <= triangle_rom(2741);
     when "101010110110" => data <= triangle_rom(2742);
     when "101010110111" => data <= triangle_rom(2743);
     when "101010111000" => data <= triangle_rom(2744);
     when "101010111001" => data <= triangle_rom(2745);
     when "101010111010" => data <= triangle_rom(2746);
     when "101010111011" => data <= triangle_rom(2747);
     when "101010111100" => data <= triangle_rom(2748);
     when "101010111101" => data <= triangle_rom(2749);
     when "101010111110" => data <= triangle_rom(2750);
     when "101010111111" => data <= triangle_rom(2751);
     when "101011000000" => data <= triangle_rom(2752);
     when "101011000001" => data <= triangle_rom(2753);
     when "101011000010" => data <= triangle_rom(2754);
     when "101011000011" => data <= triangle_rom(2755);
     when "101011000100" => data <= triangle_rom(2756);
     when "101011000101" => data <= triangle_rom(2757);
     when "101011000110" => data <= triangle_rom(2758);
     when "101011000111" => data <= triangle_rom(2759);
     when "101011001000" => data <= triangle_rom(2760);
     when "101011001001" => data <= triangle_rom(2761);
     when "101011001010" => data <= triangle_rom(2762);
     when "101011001011" => data <= triangle_rom(2763);
     when "101011001100" => data <= triangle_rom(2764);
     when "101011001101" => data <= triangle_rom(2765);
     when "101011001110" => data <= triangle_rom(2766);
     when "101011001111" => data <= triangle_rom(2767);
     when "101011010000" => data <= triangle_rom(2768);
     when "101011010001" => data <= triangle_rom(2769);
     when "101011010010" => data <= triangle_rom(2770);
     when "101011010011" => data <= triangle_rom(2771);
     when "101011010100" => data <= triangle_rom(2772);
     when "101011010101" => data <= triangle_rom(2773);
     when "101011010110" => data <= triangle_rom(2774);
     when "101011010111" => data <= triangle_rom(2775);
     when "101011011000" => data <= triangle_rom(2776);
     when "101011011001" => data <= triangle_rom(2777);
     when "101011011010" => data <= triangle_rom(2778);
     when "101011011011" => data <= triangle_rom(2779);
     when "101011011100" => data <= triangle_rom(2780);
     when "101011011101" => data <= triangle_rom(2781);
     when "101011011110" => data <= triangle_rom(2782);
     when "101011011111" => data <= triangle_rom(2783);
     when "101011100000" => data <= triangle_rom(2784);
     when "101011100001" => data <= triangle_rom(2785);
     when "101011100010" => data <= triangle_rom(2786);
     when "101011100011" => data <= triangle_rom(2787);
     when "101011100100" => data <= triangle_rom(2788);
     when "101011100101" => data <= triangle_rom(2789);
     when "101011100110" => data <= triangle_rom(2790);
     when "101011100111" => data <= triangle_rom(2791);
     when "101011101000" => data <= triangle_rom(2792);
     when "101011101001" => data <= triangle_rom(2793);
     when "101011101010" => data <= triangle_rom(2794);
     when "101011101011" => data <= triangle_rom(2795);
     when "101011101100" => data <= triangle_rom(2796);
     when "101011101101" => data <= triangle_rom(2797);
     when "101011101110" => data <= triangle_rom(2798);
     when "101011101111" => data <= triangle_rom(2799);
     when "101011110000" => data <= triangle_rom(2800);
     when "101011110001" => data <= triangle_rom(2801);
     when "101011110010" => data <= triangle_rom(2802);
     when "101011110011" => data <= triangle_rom(2803);
     when "101011110100" => data <= triangle_rom(2804);
     when "101011110101" => data <= triangle_rom(2805);
     when "101011110110" => data <= triangle_rom(2806);
     when "101011110111" => data <= triangle_rom(2807);
     when "101011111000" => data <= triangle_rom(2808);
     when "101011111001" => data <= triangle_rom(2809);
     when "101011111010" => data <= triangle_rom(2810);
     when "101011111011" => data <= triangle_rom(2811);
     when "101011111100" => data <= triangle_rom(2812);
     when "101011111101" => data <= triangle_rom(2813);
     when "101011111110" => data <= triangle_rom(2814);
     when "101011111111" => data <= triangle_rom(2815);
     when "101100000000" => data <= triangle_rom(2816);
     when "101100000001" => data <= triangle_rom(2817);
     when "101100000010" => data <= triangle_rom(2818);
     when "101100000011" => data <= triangle_rom(2819);
     when "101100000100" => data <= triangle_rom(2820);
     when "101100000101" => data <= triangle_rom(2821);
     when "101100000110" => data <= triangle_rom(2822);
     when "101100000111" => data <= triangle_rom(2823);
     when "101100001000" => data <= triangle_rom(2824);
     when "101100001001" => data <= triangle_rom(2825);
     when "101100001010" => data <= triangle_rom(2826);
     when "101100001011" => data <= triangle_rom(2827);
     when "101100001100" => data <= triangle_rom(2828);
     when "101100001101" => data <= triangle_rom(2829);
     when "101100001110" => data <= triangle_rom(2830);
     when "101100001111" => data <= triangle_rom(2831);
     when "101100010000" => data <= triangle_rom(2832);
     when "101100010001" => data <= triangle_rom(2833);
     when "101100010010" => data <= triangle_rom(2834);
     when "101100010011" => data <= triangle_rom(2835);
     when "101100010100" => data <= triangle_rom(2836);
     when "101100010101" => data <= triangle_rom(2837);
     when "101100010110" => data <= triangle_rom(2838);
     when "101100010111" => data <= triangle_rom(2839);
     when "101100011000" => data <= triangle_rom(2840);
     when "101100011001" => data <= triangle_rom(2841);
     when "101100011010" => data <= triangle_rom(2842);
     when "101100011011" => data <= triangle_rom(2843);
     when "101100011100" => data <= triangle_rom(2844);
     when "101100011101" => data <= triangle_rom(2845);
     when "101100011110" => data <= triangle_rom(2846);
     when "101100011111" => data <= triangle_rom(2847);
     when "101100100000" => data <= triangle_rom(2848);
     when "101100100001" => data <= triangle_rom(2849);
     when "101100100010" => data <= triangle_rom(2850);
     when "101100100011" => data <= triangle_rom(2851);
     when "101100100100" => data <= triangle_rom(2852);
     when "101100100101" => data <= triangle_rom(2853);
     when "101100100110" => data <= triangle_rom(2854);
     when "101100100111" => data <= triangle_rom(2855);
     when "101100101000" => data <= triangle_rom(2856);
     when "101100101001" => data <= triangle_rom(2857);
     when "101100101010" => data <= triangle_rom(2858);
     when "101100101011" => data <= triangle_rom(2859);
     when "101100101100" => data <= triangle_rom(2860);
     when "101100101101" => data <= triangle_rom(2861);
     when "101100101110" => data <= triangle_rom(2862);
     when "101100101111" => data <= triangle_rom(2863);
     when "101100110000" => data <= triangle_rom(2864);
     when "101100110001" => data <= triangle_rom(2865);
     when "101100110010" => data <= triangle_rom(2866);
     when "101100110011" => data <= triangle_rom(2867);
     when "101100110100" => data <= triangle_rom(2868);
     when "101100110101" => data <= triangle_rom(2869);
     when "101100110110" => data <= triangle_rom(2870);
     when "101100110111" => data <= triangle_rom(2871);
     when "101100111000" => data <= triangle_rom(2872);
     when "101100111001" => data <= triangle_rom(2873);
     when "101100111010" => data <= triangle_rom(2874);
     when "101100111011" => data <= triangle_rom(2875);
     when "101100111100" => data <= triangle_rom(2876);
     when "101100111101" => data <= triangle_rom(2877);
     when "101100111110" => data <= triangle_rom(2878);
     when "101100111111" => data <= triangle_rom(2879);
     when "101101000000" => data <= triangle_rom(2880);
     when "101101000001" => data <= triangle_rom(2881);
     when "101101000010" => data <= triangle_rom(2882);
     when "101101000011" => data <= triangle_rom(2883);
     when "101101000100" => data <= triangle_rom(2884);
     when "101101000101" => data <= triangle_rom(2885);
     when "101101000110" => data <= triangle_rom(2886);
     when "101101000111" => data <= triangle_rom(2887);
     when "101101001000" => data <= triangle_rom(2888);
     when "101101001001" => data <= triangle_rom(2889);
     when "101101001010" => data <= triangle_rom(2890);
     when "101101001011" => data <= triangle_rom(2891);
     when "101101001100" => data <= triangle_rom(2892);
     when "101101001101" => data <= triangle_rom(2893);
     when "101101001110" => data <= triangle_rom(2894);
     when "101101001111" => data <= triangle_rom(2895);
     when "101101010000" => data <= triangle_rom(2896);
     when "101101010001" => data <= triangle_rom(2897);
     when "101101010010" => data <= triangle_rom(2898);
     when "101101010011" => data <= triangle_rom(2899);
     when "101101010100" => data <= triangle_rom(2900);
     when "101101010101" => data <= triangle_rom(2901);
     when "101101010110" => data <= triangle_rom(2902);
     when "101101010111" => data <= triangle_rom(2903);
     when "101101011000" => data <= triangle_rom(2904);
     when "101101011001" => data <= triangle_rom(2905);
     when "101101011010" => data <= triangle_rom(2906);
     when "101101011011" => data <= triangle_rom(2907);
     when "101101011100" => data <= triangle_rom(2908);
     when "101101011101" => data <= triangle_rom(2909);
     when "101101011110" => data <= triangle_rom(2910);
     when "101101011111" => data <= triangle_rom(2911);
     when "101101100000" => data <= triangle_rom(2912);
     when "101101100001" => data <= triangle_rom(2913);
     when "101101100010" => data <= triangle_rom(2914);
     when "101101100011" => data <= triangle_rom(2915);
     when "101101100100" => data <= triangle_rom(2916);
     when "101101100101" => data <= triangle_rom(2917);
     when "101101100110" => data <= triangle_rom(2918);
     when "101101100111" => data <= triangle_rom(2919);
     when "101101101000" => data <= triangle_rom(2920);
     when "101101101001" => data <= triangle_rom(2921);
     when "101101101010" => data <= triangle_rom(2922);
     when "101101101011" => data <= triangle_rom(2923);
     when "101101101100" => data <= triangle_rom(2924);
     when "101101101101" => data <= triangle_rom(2925);
     when "101101101110" => data <= triangle_rom(2926);
     when "101101101111" => data <= triangle_rom(2927);
     when "101101110000" => data <= triangle_rom(2928);
     when "101101110001" => data <= triangle_rom(2929);
     when "101101110010" => data <= triangle_rom(2930);
     when "101101110011" => data <= triangle_rom(2931);
     when "101101110100" => data <= triangle_rom(2932);
     when "101101110101" => data <= triangle_rom(2933);
     when "101101110110" => data <= triangle_rom(2934);
     when "101101110111" => data <= triangle_rom(2935);
     when "101101111000" => data <= triangle_rom(2936);
     when "101101111001" => data <= triangle_rom(2937);
     when "101101111010" => data <= triangle_rom(2938);
     when "101101111011" => data <= triangle_rom(2939);
     when "101101111100" => data <= triangle_rom(2940);
     when "101101111101" => data <= triangle_rom(2941);
     when "101101111110" => data <= triangle_rom(2942);
     when "101101111111" => data <= triangle_rom(2943);
     when "101110000000" => data <= triangle_rom(2944);
     when "101110000001" => data <= triangle_rom(2945);
     when "101110000010" => data <= triangle_rom(2946);
     when "101110000011" => data <= triangle_rom(2947);
     when "101110000100" => data <= triangle_rom(2948);
     when "101110000101" => data <= triangle_rom(2949);
     when "101110000110" => data <= triangle_rom(2950);
     when "101110000111" => data <= triangle_rom(2951);
     when "101110001000" => data <= triangle_rom(2952);
     when "101110001001" => data <= triangle_rom(2953);
     when "101110001010" => data <= triangle_rom(2954);
     when "101110001011" => data <= triangle_rom(2955);
     when "101110001100" => data <= triangle_rom(2956);
     when "101110001101" => data <= triangle_rom(2957);
     when "101110001110" => data <= triangle_rom(2958);
     when "101110001111" => data <= triangle_rom(2959);
     when "101110010000" => data <= triangle_rom(2960);
     when "101110010001" => data <= triangle_rom(2961);
     when "101110010010" => data <= triangle_rom(2962);
     when "101110010011" => data <= triangle_rom(2963);
     when "101110010100" => data <= triangle_rom(2964);
     when "101110010101" => data <= triangle_rom(2965);
     when "101110010110" => data <= triangle_rom(2966);
     when "101110010111" => data <= triangle_rom(2967);
     when "101110011000" => data <= triangle_rom(2968);
     when "101110011001" => data <= triangle_rom(2969);
     when "101110011010" => data <= triangle_rom(2970);
     when "101110011011" => data <= triangle_rom(2971);
     when "101110011100" => data <= triangle_rom(2972);
     when "101110011101" => data <= triangle_rom(2973);
     when "101110011110" => data <= triangle_rom(2974);
     when "101110011111" => data <= triangle_rom(2975);
     when "101110100000" => data <= triangle_rom(2976);
     when "101110100001" => data <= triangle_rom(2977);
     when "101110100010" => data <= triangle_rom(2978);
     when "101110100011" => data <= triangle_rom(2979);
     when "101110100100" => data <= triangle_rom(2980);
     when "101110100101" => data <= triangle_rom(2981);
     when "101110100110" => data <= triangle_rom(2982);
     when "101110100111" => data <= triangle_rom(2983);
     when "101110101000" => data <= triangle_rom(2984);
     when "101110101001" => data <= triangle_rom(2985);
     when "101110101010" => data <= triangle_rom(2986);
     when "101110101011" => data <= triangle_rom(2987);
     when "101110101100" => data <= triangle_rom(2988);
     when "101110101101" => data <= triangle_rom(2989);
     when "101110101110" => data <= triangle_rom(2990);
     when "101110101111" => data <= triangle_rom(2991);
     when "101110110000" => data <= triangle_rom(2992);
     when "101110110001" => data <= triangle_rom(2993);
     when "101110110010" => data <= triangle_rom(2994);
     when "101110110011" => data <= triangle_rom(2995);
     when "101110110100" => data <= triangle_rom(2996);
     when "101110110101" => data <= triangle_rom(2997);
     when "101110110110" => data <= triangle_rom(2998);
     when "101110110111" => data <= triangle_rom(2999);
     when "101110111000" => data <= triangle_rom(3000);
     when "101110111001" => data <= triangle_rom(3001);
     when "101110111010" => data <= triangle_rom(3002);
     when "101110111011" => data <= triangle_rom(3003);
     when "101110111100" => data <= triangle_rom(3004);
     when "101110111101" => data <= triangle_rom(3005);
     when "101110111110" => data <= triangle_rom(3006);
     when "101110111111" => data <= triangle_rom(3007);
     when "101111000000" => data <= triangle_rom(3008);
     when "101111000001" => data <= triangle_rom(3009);
     when "101111000010" => data <= triangle_rom(3010);
     when "101111000011" => data <= triangle_rom(3011);
     when "101111000100" => data <= triangle_rom(3012);
     when "101111000101" => data <= triangle_rom(3013);
     when "101111000110" => data <= triangle_rom(3014);
     when "101111000111" => data <= triangle_rom(3015);
     when "101111001000" => data <= triangle_rom(3016);
     when "101111001001" => data <= triangle_rom(3017);
     when "101111001010" => data <= triangle_rom(3018);
     when "101111001011" => data <= triangle_rom(3019);
     when "101111001100" => data <= triangle_rom(3020);
     when "101111001101" => data <= triangle_rom(3021);
     when "101111001110" => data <= triangle_rom(3022);
     when "101111001111" => data <= triangle_rom(3023);
     when "101111010000" => data <= triangle_rom(3024);
     when "101111010001" => data <= triangle_rom(3025);
     when "101111010010" => data <= triangle_rom(3026);
     when "101111010011" => data <= triangle_rom(3027);
     when "101111010100" => data <= triangle_rom(3028);
     when "101111010101" => data <= triangle_rom(3029);
     when "101111010110" => data <= triangle_rom(3030);
     when "101111010111" => data <= triangle_rom(3031);
     when "101111011000" => data <= triangle_rom(3032);
     when "101111011001" => data <= triangle_rom(3033);
     when "101111011010" => data <= triangle_rom(3034);
     when "101111011011" => data <= triangle_rom(3035);
     when "101111011100" => data <= triangle_rom(3036);
     when "101111011101" => data <= triangle_rom(3037);
     when "101111011110" => data <= triangle_rom(3038);
     when "101111011111" => data <= triangle_rom(3039);
     when "101111100000" => data <= triangle_rom(3040);
     when "101111100001" => data <= triangle_rom(3041);
     when "101111100010" => data <= triangle_rom(3042);
     when "101111100011" => data <= triangle_rom(3043);
     when "101111100100" => data <= triangle_rom(3044);
     when "101111100101" => data <= triangle_rom(3045);
     when "101111100110" => data <= triangle_rom(3046);
     when "101111100111" => data <= triangle_rom(3047);
     when "101111101000" => data <= triangle_rom(3048);
     when "101111101001" => data <= triangle_rom(3049);
     when "101111101010" => data <= triangle_rom(3050);
     when "101111101011" => data <= triangle_rom(3051);
     when "101111101100" => data <= triangle_rom(3052);
     when "101111101101" => data <= triangle_rom(3053);
     when "101111101110" => data <= triangle_rom(3054);
     when "101111101111" => data <= triangle_rom(3055);
     when "101111110000" => data <= triangle_rom(3056);
     when "101111110001" => data <= triangle_rom(3057);
     when "101111110010" => data <= triangle_rom(3058);
     when "101111110011" => data <= triangle_rom(3059);
     when "101111110100" => data <= triangle_rom(3060);
     when "101111110101" => data <= triangle_rom(3061);
     when "101111110110" => data <= triangle_rom(3062);
     when "101111110111" => data <= triangle_rom(3063);
     when "101111111000" => data <= triangle_rom(3064);
     when "101111111001" => data <= triangle_rom(3065);
     when "101111111010" => data <= triangle_rom(3066);
     when "101111111011" => data <= triangle_rom(3067);
     when "101111111100" => data <= triangle_rom(3068);
     when "101111111101" => data <= triangle_rom(3069);
     when "101111111110" => data <= triangle_rom(3070);
     when "101111111111" => data <= triangle_rom(3071);
     when "110000000000" => data <= triangle_rom(3072);
     when "110000000001" => data <= triangle_rom(3073);
     when "110000000010" => data <= triangle_rom(3074);
     when "110000000011" => data <= triangle_rom(3075);
     when "110000000100" => data <= triangle_rom(3076);
     when "110000000101" => data <= triangle_rom(3077);
     when "110000000110" => data <= triangle_rom(3078);
     when "110000000111" => data <= triangle_rom(3079);
     when "110000001000" => data <= triangle_rom(3080);
     when "110000001001" => data <= triangle_rom(3081);
     when "110000001010" => data <= triangle_rom(3082);
     when "110000001011" => data <= triangle_rom(3083);
     when "110000001100" => data <= triangle_rom(3084);
     when "110000001101" => data <= triangle_rom(3085);
     when "110000001110" => data <= triangle_rom(3086);
     when "110000001111" => data <= triangle_rom(3087);
     when "110000010000" => data <= triangle_rom(3088);
     when "110000010001" => data <= triangle_rom(3089);
     when "110000010010" => data <= triangle_rom(3090);
     when "110000010011" => data <= triangle_rom(3091);
     when "110000010100" => data <= triangle_rom(3092);
     when "110000010101" => data <= triangle_rom(3093);
     when "110000010110" => data <= triangle_rom(3094);
     when "110000010111" => data <= triangle_rom(3095);
     when "110000011000" => data <= triangle_rom(3096);
     when "110000011001" => data <= triangle_rom(3097);
     when "110000011010" => data <= triangle_rom(3098);
     when "110000011011" => data <= triangle_rom(3099);
     when "110000011100" => data <= triangle_rom(3100);
     when "110000011101" => data <= triangle_rom(3101);
     when "110000011110" => data <= triangle_rom(3102);
     when "110000011111" => data <= triangle_rom(3103);
     when "110000100000" => data <= triangle_rom(3104);
     when "110000100001" => data <= triangle_rom(3105);
     when "110000100010" => data <= triangle_rom(3106);
     when "110000100011" => data <= triangle_rom(3107);
     when "110000100100" => data <= triangle_rom(3108);
     when "110000100101" => data <= triangle_rom(3109);
     when "110000100110" => data <= triangle_rom(3110);
     when "110000100111" => data <= triangle_rom(3111);
     when "110000101000" => data <= triangle_rom(3112);
     when "110000101001" => data <= triangle_rom(3113);
     when "110000101010" => data <= triangle_rom(3114);
     when "110000101011" => data <= triangle_rom(3115);
     when "110000101100" => data <= triangle_rom(3116);
     when "110000101101" => data <= triangle_rom(3117);
     when "110000101110" => data <= triangle_rom(3118);
     when "110000101111" => data <= triangle_rom(3119);
     when "110000110000" => data <= triangle_rom(3120);
     when "110000110001" => data <= triangle_rom(3121);
     when "110000110010" => data <= triangle_rom(3122);
     when "110000110011" => data <= triangle_rom(3123);
     when "110000110100" => data <= triangle_rom(3124);
     when "110000110101" => data <= triangle_rom(3125);
     when "110000110110" => data <= triangle_rom(3126);
     when "110000110111" => data <= triangle_rom(3127);
     when "110000111000" => data <= triangle_rom(3128);
     when "110000111001" => data <= triangle_rom(3129);
     when "110000111010" => data <= triangle_rom(3130);
     when "110000111011" => data <= triangle_rom(3131);
     when "110000111100" => data <= triangle_rom(3132);
     when "110000111101" => data <= triangle_rom(3133);
     when "110000111110" => data <= triangle_rom(3134);
     when "110000111111" => data <= triangle_rom(3135);
     when "110001000000" => data <= triangle_rom(3136);
     when "110001000001" => data <= triangle_rom(3137);
     when "110001000010" => data <= triangle_rom(3138);
     when "110001000011" => data <= triangle_rom(3139);
     when "110001000100" => data <= triangle_rom(3140);
     when "110001000101" => data <= triangle_rom(3141);
     when "110001000110" => data <= triangle_rom(3142);
     when "110001000111" => data <= triangle_rom(3143);
     when "110001001000" => data <= triangle_rom(3144);
     when "110001001001" => data <= triangle_rom(3145);
     when "110001001010" => data <= triangle_rom(3146);
     when "110001001011" => data <= triangle_rom(3147);
     when "110001001100" => data <= triangle_rom(3148);
     when "110001001101" => data <= triangle_rom(3149);
     when "110001001110" => data <= triangle_rom(3150);
     when "110001001111" => data <= triangle_rom(3151);
     when "110001010000" => data <= triangle_rom(3152);
     when "110001010001" => data <= triangle_rom(3153);
     when "110001010010" => data <= triangle_rom(3154);
     when "110001010011" => data <= triangle_rom(3155);
     when "110001010100" => data <= triangle_rom(3156);
     when "110001010101" => data <= triangle_rom(3157);
     when "110001010110" => data <= triangle_rom(3158);
     when "110001010111" => data <= triangle_rom(3159);
     when "110001011000" => data <= triangle_rom(3160);
     when "110001011001" => data <= triangle_rom(3161);
     when "110001011010" => data <= triangle_rom(3162);
     when "110001011011" => data <= triangle_rom(3163);
     when "110001011100" => data <= triangle_rom(3164);
     when "110001011101" => data <= triangle_rom(3165);
     when "110001011110" => data <= triangle_rom(3166);
     when "110001011111" => data <= triangle_rom(3167);
     when "110001100000" => data <= triangle_rom(3168);
     when "110001100001" => data <= triangle_rom(3169);
     when "110001100010" => data <= triangle_rom(3170);
     when "110001100011" => data <= triangle_rom(3171);
     when "110001100100" => data <= triangle_rom(3172);
     when "110001100101" => data <= triangle_rom(3173);
     when "110001100110" => data <= triangle_rom(3174);
     when "110001100111" => data <= triangle_rom(3175);
     when "110001101000" => data <= triangle_rom(3176);
     when "110001101001" => data <= triangle_rom(3177);
     when "110001101010" => data <= triangle_rom(3178);
     when "110001101011" => data <= triangle_rom(3179);
     when "110001101100" => data <= triangle_rom(3180);
     when "110001101101" => data <= triangle_rom(3181);
     when "110001101110" => data <= triangle_rom(3182);
     when "110001101111" => data <= triangle_rom(3183);
     when "110001110000" => data <= triangle_rom(3184);
     when "110001110001" => data <= triangle_rom(3185);
     when "110001110010" => data <= triangle_rom(3186);
     when "110001110011" => data <= triangle_rom(3187);
     when "110001110100" => data <= triangle_rom(3188);
     when "110001110101" => data <= triangle_rom(3189);
     when "110001110110" => data <= triangle_rom(3190);
     when "110001110111" => data <= triangle_rom(3191);
     when "110001111000" => data <= triangle_rom(3192);
     when "110001111001" => data <= triangle_rom(3193);
     when "110001111010" => data <= triangle_rom(3194);
     when "110001111011" => data <= triangle_rom(3195);
     when "110001111100" => data <= triangle_rom(3196);
     when "110001111101" => data <= triangle_rom(3197);
     when "110001111110" => data <= triangle_rom(3198);
     when "110001111111" => data <= triangle_rom(3199);
     when "110010000000" => data <= triangle_rom(3200);
     when "110010000001" => data <= triangle_rom(3201);
     when "110010000010" => data <= triangle_rom(3202);
     when "110010000011" => data <= triangle_rom(3203);
     when "110010000100" => data <= triangle_rom(3204);
     when "110010000101" => data <= triangle_rom(3205);
     when "110010000110" => data <= triangle_rom(3206);
     when "110010000111" => data <= triangle_rom(3207);
     when "110010001000" => data <= triangle_rom(3208);
     when "110010001001" => data <= triangle_rom(3209);
     when "110010001010" => data <= triangle_rom(3210);
     when "110010001011" => data <= triangle_rom(3211);
     when "110010001100" => data <= triangle_rom(3212);
     when "110010001101" => data <= triangle_rom(3213);
     when "110010001110" => data <= triangle_rom(3214);
     when "110010001111" => data <= triangle_rom(3215);
     when "110010010000" => data <= triangle_rom(3216);
     when "110010010001" => data <= triangle_rom(3217);
     when "110010010010" => data <= triangle_rom(3218);
     when "110010010011" => data <= triangle_rom(3219);
     when "110010010100" => data <= triangle_rom(3220);
     when "110010010101" => data <= triangle_rom(3221);
     when "110010010110" => data <= triangle_rom(3222);
     when "110010010111" => data <= triangle_rom(3223);
     when "110010011000" => data <= triangle_rom(3224);
     when "110010011001" => data <= triangle_rom(3225);
     when "110010011010" => data <= triangle_rom(3226);
     when "110010011011" => data <= triangle_rom(3227);
     when "110010011100" => data <= triangle_rom(3228);
     when "110010011101" => data <= triangle_rom(3229);
     when "110010011110" => data <= triangle_rom(3230);
     when "110010011111" => data <= triangle_rom(3231);
     when "110010100000" => data <= triangle_rom(3232);
     when "110010100001" => data <= triangle_rom(3233);
     when "110010100010" => data <= triangle_rom(3234);
     when "110010100011" => data <= triangle_rom(3235);
     when "110010100100" => data <= triangle_rom(3236);
     when "110010100101" => data <= triangle_rom(3237);
     when "110010100110" => data <= triangle_rom(3238);
     when "110010100111" => data <= triangle_rom(3239);
     when "110010101000" => data <= triangle_rom(3240);
     when "110010101001" => data <= triangle_rom(3241);
     when "110010101010" => data <= triangle_rom(3242);
     when "110010101011" => data <= triangle_rom(3243);
     when "110010101100" => data <= triangle_rom(3244);
     when "110010101101" => data <= triangle_rom(3245);
     when "110010101110" => data <= triangle_rom(3246);
     when "110010101111" => data <= triangle_rom(3247);
     when "110010110000" => data <= triangle_rom(3248);
     when "110010110001" => data <= triangle_rom(3249);
     when "110010110010" => data <= triangle_rom(3250);
     when "110010110011" => data <= triangle_rom(3251);
     when "110010110100" => data <= triangle_rom(3252);
     when "110010110101" => data <= triangle_rom(3253);
     when "110010110110" => data <= triangle_rom(3254);
     when "110010110111" => data <= triangle_rom(3255);
     when "110010111000" => data <= triangle_rom(3256);
     when "110010111001" => data <= triangle_rom(3257);
     when "110010111010" => data <= triangle_rom(3258);
     when "110010111011" => data <= triangle_rom(3259);
     when "110010111100" => data <= triangle_rom(3260);
     when "110010111101" => data <= triangle_rom(3261);
     when "110010111110" => data <= triangle_rom(3262);
     when "110010111111" => data <= triangle_rom(3263);
     when "110011000000" => data <= triangle_rom(3264);
     when "110011000001" => data <= triangle_rom(3265);
     when "110011000010" => data <= triangle_rom(3266);
     when "110011000011" => data <= triangle_rom(3267);
     when "110011000100" => data <= triangle_rom(3268);
     when "110011000101" => data <= triangle_rom(3269);
     when "110011000110" => data <= triangle_rom(3270);
     when "110011000111" => data <= triangle_rom(3271);
     when "110011001000" => data <= triangle_rom(3272);
     when "110011001001" => data <= triangle_rom(3273);
     when "110011001010" => data <= triangle_rom(3274);
     when "110011001011" => data <= triangle_rom(3275);
     when "110011001100" => data <= triangle_rom(3276);
     when "110011001101" => data <= triangle_rom(3277);
     when "110011001110" => data <= triangle_rom(3278);
     when "110011001111" => data <= triangle_rom(3279);
     when "110011010000" => data <= triangle_rom(3280);
     when "110011010001" => data <= triangle_rom(3281);
     when "110011010010" => data <= triangle_rom(3282);
     when "110011010011" => data <= triangle_rom(3283);
     when "110011010100" => data <= triangle_rom(3284);
     when "110011010101" => data <= triangle_rom(3285);
     when "110011010110" => data <= triangle_rom(3286);
     when "110011010111" => data <= triangle_rom(3287);
     when "110011011000" => data <= triangle_rom(3288);
     when "110011011001" => data <= triangle_rom(3289);
     when "110011011010" => data <= triangle_rom(3290);
     when "110011011011" => data <= triangle_rom(3291);
     when "110011011100" => data <= triangle_rom(3292);
     when "110011011101" => data <= triangle_rom(3293);
     when "110011011110" => data <= triangle_rom(3294);
     when "110011011111" => data <= triangle_rom(3295);
     when "110011100000" => data <= triangle_rom(3296);
     when "110011100001" => data <= triangle_rom(3297);
     when "110011100010" => data <= triangle_rom(3298);
     when "110011100011" => data <= triangle_rom(3299);
     when "110011100100" => data <= triangle_rom(3300);
     when "110011100101" => data <= triangle_rom(3301);
     when "110011100110" => data <= triangle_rom(3302);
     when "110011100111" => data <= triangle_rom(3303);
     when "110011101000" => data <= triangle_rom(3304);
     when "110011101001" => data <= triangle_rom(3305);
     when "110011101010" => data <= triangle_rom(3306);
     when "110011101011" => data <= triangle_rom(3307);
     when "110011101100" => data <= triangle_rom(3308);
     when "110011101101" => data <= triangle_rom(3309);
     when "110011101110" => data <= triangle_rom(3310);
     when "110011101111" => data <= triangle_rom(3311);
     when "110011110000" => data <= triangle_rom(3312);
     when "110011110001" => data <= triangle_rom(3313);
     when "110011110010" => data <= triangle_rom(3314);
     when "110011110011" => data <= triangle_rom(3315);
     when "110011110100" => data <= triangle_rom(3316);
     when "110011110101" => data <= triangle_rom(3317);
     when "110011110110" => data <= triangle_rom(3318);
     when "110011110111" => data <= triangle_rom(3319);
     when "110011111000" => data <= triangle_rom(3320);
     when "110011111001" => data <= triangle_rom(3321);
     when "110011111010" => data <= triangle_rom(3322);
     when "110011111011" => data <= triangle_rom(3323);
     when "110011111100" => data <= triangle_rom(3324);
     when "110011111101" => data <= triangle_rom(3325);
     when "110011111110" => data <= triangle_rom(3326);
     when "110011111111" => data <= triangle_rom(3327);
     when "110100000000" => data <= triangle_rom(3328);
     when "110100000001" => data <= triangle_rom(3329);
     when "110100000010" => data <= triangle_rom(3330);
     when "110100000011" => data <= triangle_rom(3331);
     when "110100000100" => data <= triangle_rom(3332);
     when "110100000101" => data <= triangle_rom(3333);
     when "110100000110" => data <= triangle_rom(3334);
     when "110100000111" => data <= triangle_rom(3335);
     when "110100001000" => data <= triangle_rom(3336);
     when "110100001001" => data <= triangle_rom(3337);
     when "110100001010" => data <= triangle_rom(3338);
     when "110100001011" => data <= triangle_rom(3339);
     when "110100001100" => data <= triangle_rom(3340);
     when "110100001101" => data <= triangle_rom(3341);
     when "110100001110" => data <= triangle_rom(3342);
     when "110100001111" => data <= triangle_rom(3343);
     when "110100010000" => data <= triangle_rom(3344);
     when "110100010001" => data <= triangle_rom(3345);
     when "110100010010" => data <= triangle_rom(3346);
     when "110100010011" => data <= triangle_rom(3347);
     when "110100010100" => data <= triangle_rom(3348);
     when "110100010101" => data <= triangle_rom(3349);
     when "110100010110" => data <= triangle_rom(3350);
     when "110100010111" => data <= triangle_rom(3351);
     when "110100011000" => data <= triangle_rom(3352);
     when "110100011001" => data <= triangle_rom(3353);
     when "110100011010" => data <= triangle_rom(3354);
     when "110100011011" => data <= triangle_rom(3355);
     when "110100011100" => data <= triangle_rom(3356);
     when "110100011101" => data <= triangle_rom(3357);
     when "110100011110" => data <= triangle_rom(3358);
     when "110100011111" => data <= triangle_rom(3359);
     when "110100100000" => data <= triangle_rom(3360);
     when "110100100001" => data <= triangle_rom(3361);
     when "110100100010" => data <= triangle_rom(3362);
     when "110100100011" => data <= triangle_rom(3363);
     when "110100100100" => data <= triangle_rom(3364);
     when "110100100101" => data <= triangle_rom(3365);
     when "110100100110" => data <= triangle_rom(3366);
     when "110100100111" => data <= triangle_rom(3367);
     when "110100101000" => data <= triangle_rom(3368);
     when "110100101001" => data <= triangle_rom(3369);
     when "110100101010" => data <= triangle_rom(3370);
     when "110100101011" => data <= triangle_rom(3371);
     when "110100101100" => data <= triangle_rom(3372);
     when "110100101101" => data <= triangle_rom(3373);
     when "110100101110" => data <= triangle_rom(3374);
     when "110100101111" => data <= triangle_rom(3375);
     when "110100110000" => data <= triangle_rom(3376);
     when "110100110001" => data <= triangle_rom(3377);
     when "110100110010" => data <= triangle_rom(3378);
     when "110100110011" => data <= triangle_rom(3379);
     when "110100110100" => data <= triangle_rom(3380);
     when "110100110101" => data <= triangle_rom(3381);
     when "110100110110" => data <= triangle_rom(3382);
     when "110100110111" => data <= triangle_rom(3383);
     when "110100111000" => data <= triangle_rom(3384);
     when "110100111001" => data <= triangle_rom(3385);
     when "110100111010" => data <= triangle_rom(3386);
     when "110100111011" => data <= triangle_rom(3387);
     when "110100111100" => data <= triangle_rom(3388);
     when "110100111101" => data <= triangle_rom(3389);
     when "110100111110" => data <= triangle_rom(3390);
     when "110100111111" => data <= triangle_rom(3391);
     when "110101000000" => data <= triangle_rom(3392);
     when "110101000001" => data <= triangle_rom(3393);
     when "110101000010" => data <= triangle_rom(3394);
     when "110101000011" => data <= triangle_rom(3395);
     when "110101000100" => data <= triangle_rom(3396);
     when "110101000101" => data <= triangle_rom(3397);
     when "110101000110" => data <= triangle_rom(3398);
     when "110101000111" => data <= triangle_rom(3399);
     when "110101001000" => data <= triangle_rom(3400);
     when "110101001001" => data <= triangle_rom(3401);
     when "110101001010" => data <= triangle_rom(3402);
     when "110101001011" => data <= triangle_rom(3403);
     when "110101001100" => data <= triangle_rom(3404);
     when "110101001101" => data <= triangle_rom(3405);
     when "110101001110" => data <= triangle_rom(3406);
     when "110101001111" => data <= triangle_rom(3407);
     when "110101010000" => data <= triangle_rom(3408);
     when "110101010001" => data <= triangle_rom(3409);
     when "110101010010" => data <= triangle_rom(3410);
     when "110101010011" => data <= triangle_rom(3411);
     when "110101010100" => data <= triangle_rom(3412);
     when "110101010101" => data <= triangle_rom(3413);
     when "110101010110" => data <= triangle_rom(3414);
     when "110101010111" => data <= triangle_rom(3415);
     when "110101011000" => data <= triangle_rom(3416);
     when "110101011001" => data <= triangle_rom(3417);
     when "110101011010" => data <= triangle_rom(3418);
     when "110101011011" => data <= triangle_rom(3419);
     when "110101011100" => data <= triangle_rom(3420);
     when "110101011101" => data <= triangle_rom(3421);
     when "110101011110" => data <= triangle_rom(3422);
     when "110101011111" => data <= triangle_rom(3423);
     when "110101100000" => data <= triangle_rom(3424);
     when "110101100001" => data <= triangle_rom(3425);
     when "110101100010" => data <= triangle_rom(3426);
     when "110101100011" => data <= triangle_rom(3427);
     when "110101100100" => data <= triangle_rom(3428);
     when "110101100101" => data <= triangle_rom(3429);
     when "110101100110" => data <= triangle_rom(3430);
     when "110101100111" => data <= triangle_rom(3431);
     when "110101101000" => data <= triangle_rom(3432);
     when "110101101001" => data <= triangle_rom(3433);
     when "110101101010" => data <= triangle_rom(3434);
     when "110101101011" => data <= triangle_rom(3435);
     when "110101101100" => data <= triangle_rom(3436);
     when "110101101101" => data <= triangle_rom(3437);
     when "110101101110" => data <= triangle_rom(3438);
     when "110101101111" => data <= triangle_rom(3439);
     when "110101110000" => data <= triangle_rom(3440);
     when "110101110001" => data <= triangle_rom(3441);
     when "110101110010" => data <= triangle_rom(3442);
     when "110101110011" => data <= triangle_rom(3443);
     when "110101110100" => data <= triangle_rom(3444);
     when "110101110101" => data <= triangle_rom(3445);
     when "110101110110" => data <= triangle_rom(3446);
     when "110101110111" => data <= triangle_rom(3447);
     when "110101111000" => data <= triangle_rom(3448);
     when "110101111001" => data <= triangle_rom(3449);
     when "110101111010" => data <= triangle_rom(3450);
     when "110101111011" => data <= triangle_rom(3451);
     when "110101111100" => data <= triangle_rom(3452);
     when "110101111101" => data <= triangle_rom(3453);
     when "110101111110" => data <= triangle_rom(3454);
     when "110101111111" => data <= triangle_rom(3455);
     when "110110000000" => data <= triangle_rom(3456);
     when "110110000001" => data <= triangle_rom(3457);
     when "110110000010" => data <= triangle_rom(3458);
     when "110110000011" => data <= triangle_rom(3459);
     when "110110000100" => data <= triangle_rom(3460);
     when "110110000101" => data <= triangle_rom(3461);
     when "110110000110" => data <= triangle_rom(3462);
     when "110110000111" => data <= triangle_rom(3463);
     when "110110001000" => data <= triangle_rom(3464);
     when "110110001001" => data <= triangle_rom(3465);
     when "110110001010" => data <= triangle_rom(3466);
     when "110110001011" => data <= triangle_rom(3467);
     when "110110001100" => data <= triangle_rom(3468);
     when "110110001101" => data <= triangle_rom(3469);
     when "110110001110" => data <= triangle_rom(3470);
     when "110110001111" => data <= triangle_rom(3471);
     when "110110010000" => data <= triangle_rom(3472);
     when "110110010001" => data <= triangle_rom(3473);
     when "110110010010" => data <= triangle_rom(3474);
     when "110110010011" => data <= triangle_rom(3475);
     when "110110010100" => data <= triangle_rom(3476);
     when "110110010101" => data <= triangle_rom(3477);
     when "110110010110" => data <= triangle_rom(3478);
     when "110110010111" => data <= triangle_rom(3479);
     when "110110011000" => data <= triangle_rom(3480);
     when "110110011001" => data <= triangle_rom(3481);
     when "110110011010" => data <= triangle_rom(3482);
     when "110110011011" => data <= triangle_rom(3483);
     when "110110011100" => data <= triangle_rom(3484);
     when "110110011101" => data <= triangle_rom(3485);
     when "110110011110" => data <= triangle_rom(3486);
     when "110110011111" => data <= triangle_rom(3487);
     when "110110100000" => data <= triangle_rom(3488);
     when "110110100001" => data <= triangle_rom(3489);
     when "110110100010" => data <= triangle_rom(3490);
     when "110110100011" => data <= triangle_rom(3491);
     when "110110100100" => data <= triangle_rom(3492);
     when "110110100101" => data <= triangle_rom(3493);
     when "110110100110" => data <= triangle_rom(3494);
     when "110110100111" => data <= triangle_rom(3495);
     when "110110101000" => data <= triangle_rom(3496);
     when "110110101001" => data <= triangle_rom(3497);
     when "110110101010" => data <= triangle_rom(3498);
     when "110110101011" => data <= triangle_rom(3499);
     when "110110101100" => data <= triangle_rom(3500);
     when "110110101101" => data <= triangle_rom(3501);
     when "110110101110" => data <= triangle_rom(3502);
     when "110110101111" => data <= triangle_rom(3503);
     when "110110110000" => data <= triangle_rom(3504);
     when "110110110001" => data <= triangle_rom(3505);
     when "110110110010" => data <= triangle_rom(3506);
     when "110110110011" => data <= triangle_rom(3507);
     when "110110110100" => data <= triangle_rom(3508);
     when "110110110101" => data <= triangle_rom(3509);
     when "110110110110" => data <= triangle_rom(3510);
     when "110110110111" => data <= triangle_rom(3511);
     when "110110111000" => data <= triangle_rom(3512);
     when "110110111001" => data <= triangle_rom(3513);
     when "110110111010" => data <= triangle_rom(3514);
     when "110110111011" => data <= triangle_rom(3515);
     when "110110111100" => data <= triangle_rom(3516);
     when "110110111101" => data <= triangle_rom(3517);
     when "110110111110" => data <= triangle_rom(3518);
     when "110110111111" => data <= triangle_rom(3519);
     when "110111000000" => data <= triangle_rom(3520);
     when "110111000001" => data <= triangle_rom(3521);
     when "110111000010" => data <= triangle_rom(3522);
     when "110111000011" => data <= triangle_rom(3523);
     when "110111000100" => data <= triangle_rom(3524);
     when "110111000101" => data <= triangle_rom(3525);
     when "110111000110" => data <= triangle_rom(3526);
     when "110111000111" => data <= triangle_rom(3527);
     when "110111001000" => data <= triangle_rom(3528);
     when "110111001001" => data <= triangle_rom(3529);
     when "110111001010" => data <= triangle_rom(3530);
     when "110111001011" => data <= triangle_rom(3531);
     when "110111001100" => data <= triangle_rom(3532);
     when "110111001101" => data <= triangle_rom(3533);
     when "110111001110" => data <= triangle_rom(3534);
     when "110111001111" => data <= triangle_rom(3535);
     when "110111010000" => data <= triangle_rom(3536);
     when "110111010001" => data <= triangle_rom(3537);
     when "110111010010" => data <= triangle_rom(3538);
     when "110111010011" => data <= triangle_rom(3539);
     when "110111010100" => data <= triangle_rom(3540);
     when "110111010101" => data <= triangle_rom(3541);
     when "110111010110" => data <= triangle_rom(3542);
     when "110111010111" => data <= triangle_rom(3543);
     when "110111011000" => data <= triangle_rom(3544);
     when "110111011001" => data <= triangle_rom(3545);
     when "110111011010" => data <= triangle_rom(3546);
     when "110111011011" => data <= triangle_rom(3547);
     when "110111011100" => data <= triangle_rom(3548);
     when "110111011101" => data <= triangle_rom(3549);
     when "110111011110" => data <= triangle_rom(3550);
     when "110111011111" => data <= triangle_rom(3551);
     when "110111100000" => data <= triangle_rom(3552);
     when "110111100001" => data <= triangle_rom(3553);
     when "110111100010" => data <= triangle_rom(3554);
     when "110111100011" => data <= triangle_rom(3555);
     when "110111100100" => data <= triangle_rom(3556);
     when "110111100101" => data <= triangle_rom(3557);
     when "110111100110" => data <= triangle_rom(3558);
     when "110111100111" => data <= triangle_rom(3559);
     when "110111101000" => data <= triangle_rom(3560);
     when "110111101001" => data <= triangle_rom(3561);
     when "110111101010" => data <= triangle_rom(3562);
     when "110111101011" => data <= triangle_rom(3563);
     when "110111101100" => data <= triangle_rom(3564);
     when "110111101101" => data <= triangle_rom(3565);
     when "110111101110" => data <= triangle_rom(3566);
     when "110111101111" => data <= triangle_rom(3567);
     when "110111110000" => data <= triangle_rom(3568);
     when "110111110001" => data <= triangle_rom(3569);
     when "110111110010" => data <= triangle_rom(3570);
     when "110111110011" => data <= triangle_rom(3571);
     when "110111110100" => data <= triangle_rom(3572);
     when "110111110101" => data <= triangle_rom(3573);
     when "110111110110" => data <= triangle_rom(3574);
     when "110111110111" => data <= triangle_rom(3575);
     when "110111111000" => data <= triangle_rom(3576);
     when "110111111001" => data <= triangle_rom(3577);
     when "110111111010" => data <= triangle_rom(3578);
     when "110111111011" => data <= triangle_rom(3579);
     when "110111111100" => data <= triangle_rom(3580);
     when "110111111101" => data <= triangle_rom(3581);
     when "110111111110" => data <= triangle_rom(3582);
     when "110111111111" => data <= triangle_rom(3583);
     when "111000000000" => data <= triangle_rom(3584);
     when "111000000001" => data <= triangle_rom(3585);
     when "111000000010" => data <= triangle_rom(3586);
     when "111000000011" => data <= triangle_rom(3587);
     when "111000000100" => data <= triangle_rom(3588);
     when "111000000101" => data <= triangle_rom(3589);
     when "111000000110" => data <= triangle_rom(3590);
     when "111000000111" => data <= triangle_rom(3591);
     when "111000001000" => data <= triangle_rom(3592);
     when "111000001001" => data <= triangle_rom(3593);
     when "111000001010" => data <= triangle_rom(3594);
     when "111000001011" => data <= triangle_rom(3595);
     when "111000001100" => data <= triangle_rom(3596);
     when "111000001101" => data <= triangle_rom(3597);
     when "111000001110" => data <= triangle_rom(3598);
     when "111000001111" => data <= triangle_rom(3599);
     when "111000010000" => data <= triangle_rom(3600);
     when "111000010001" => data <= triangle_rom(3601);
     when "111000010010" => data <= triangle_rom(3602);
     when "111000010011" => data <= triangle_rom(3603);
     when "111000010100" => data <= triangle_rom(3604);
     when "111000010101" => data <= triangle_rom(3605);
     when "111000010110" => data <= triangle_rom(3606);
     when "111000010111" => data <= triangle_rom(3607);
     when "111000011000" => data <= triangle_rom(3608);
     when "111000011001" => data <= triangle_rom(3609);
     when "111000011010" => data <= triangle_rom(3610);
     when "111000011011" => data <= triangle_rom(3611);
     when "111000011100" => data <= triangle_rom(3612);
     when "111000011101" => data <= triangle_rom(3613);
     when "111000011110" => data <= triangle_rom(3614);
     when "111000011111" => data <= triangle_rom(3615);
     when "111000100000" => data <= triangle_rom(3616);
     when "111000100001" => data <= triangle_rom(3617);
     when "111000100010" => data <= triangle_rom(3618);
     when "111000100011" => data <= triangle_rom(3619);
     when "111000100100" => data <= triangle_rom(3620);
     when "111000100101" => data <= triangle_rom(3621);
     when "111000100110" => data <= triangle_rom(3622);
     when "111000100111" => data <= triangle_rom(3623);
     when "111000101000" => data <= triangle_rom(3624);
     when "111000101001" => data <= triangle_rom(3625);
     when "111000101010" => data <= triangle_rom(3626);
     when "111000101011" => data <= triangle_rom(3627);
     when "111000101100" => data <= triangle_rom(3628);
     when "111000101101" => data <= triangle_rom(3629);
     when "111000101110" => data <= triangle_rom(3630);
     when "111000101111" => data <= triangle_rom(3631);
     when "111000110000" => data <= triangle_rom(3632);
     when "111000110001" => data <= triangle_rom(3633);
     when "111000110010" => data <= triangle_rom(3634);
     when "111000110011" => data <= triangle_rom(3635);
     when "111000110100" => data <= triangle_rom(3636);
     when "111000110101" => data <= triangle_rom(3637);
     when "111000110110" => data <= triangle_rom(3638);
     when "111000110111" => data <= triangle_rom(3639);
     when "111000111000" => data <= triangle_rom(3640);
     when "111000111001" => data <= triangle_rom(3641);
     when "111000111010" => data <= triangle_rom(3642);
     when "111000111011" => data <= triangle_rom(3643);
     when "111000111100" => data <= triangle_rom(3644);
     when "111000111101" => data <= triangle_rom(3645);
     when "111000111110" => data <= triangle_rom(3646);
     when "111000111111" => data <= triangle_rom(3647);
     when "111001000000" => data <= triangle_rom(3648);
     when "111001000001" => data <= triangle_rom(3649);
     when "111001000010" => data <= triangle_rom(3650);
     when "111001000011" => data <= triangle_rom(3651);
     when "111001000100" => data <= triangle_rom(3652);
     when "111001000101" => data <= triangle_rom(3653);
     when "111001000110" => data <= triangle_rom(3654);
     when "111001000111" => data <= triangle_rom(3655);
     when "111001001000" => data <= triangle_rom(3656);
     when "111001001001" => data <= triangle_rom(3657);
     when "111001001010" => data <= triangle_rom(3658);
     when "111001001011" => data <= triangle_rom(3659);
     when "111001001100" => data <= triangle_rom(3660);
     when "111001001101" => data <= triangle_rom(3661);
     when "111001001110" => data <= triangle_rom(3662);
     when "111001001111" => data <= triangle_rom(3663);
     when "111001010000" => data <= triangle_rom(3664);
     when "111001010001" => data <= triangle_rom(3665);
     when "111001010010" => data <= triangle_rom(3666);
     when "111001010011" => data <= triangle_rom(3667);
     when "111001010100" => data <= triangle_rom(3668);
     when "111001010101" => data <= triangle_rom(3669);
     when "111001010110" => data <= triangle_rom(3670);
     when "111001010111" => data <= triangle_rom(3671);
     when "111001011000" => data <= triangle_rom(3672);
     when "111001011001" => data <= triangle_rom(3673);
     when "111001011010" => data <= triangle_rom(3674);
     when "111001011011" => data <= triangle_rom(3675);
     when "111001011100" => data <= triangle_rom(3676);
     when "111001011101" => data <= triangle_rom(3677);
     when "111001011110" => data <= triangle_rom(3678);
     when "111001011111" => data <= triangle_rom(3679);
     when "111001100000" => data <= triangle_rom(3680);
     when "111001100001" => data <= triangle_rom(3681);
     when "111001100010" => data <= triangle_rom(3682);
     when "111001100011" => data <= triangle_rom(3683);
     when "111001100100" => data <= triangle_rom(3684);
     when "111001100101" => data <= triangle_rom(3685);
     when "111001100110" => data <= triangle_rom(3686);
     when "111001100111" => data <= triangle_rom(3687);
     when "111001101000" => data <= triangle_rom(3688);
     when "111001101001" => data <= triangle_rom(3689);
     when "111001101010" => data <= triangle_rom(3690);
     when "111001101011" => data <= triangle_rom(3691);
     when "111001101100" => data <= triangle_rom(3692);
     when "111001101101" => data <= triangle_rom(3693);
     when "111001101110" => data <= triangle_rom(3694);
     when "111001101111" => data <= triangle_rom(3695);
     when "111001110000" => data <= triangle_rom(3696);
     when "111001110001" => data <= triangle_rom(3697);
     when "111001110010" => data <= triangle_rom(3698);
     when "111001110011" => data <= triangle_rom(3699);
     when "111001110100" => data <= triangle_rom(3700);
     when "111001110101" => data <= triangle_rom(3701);
     when "111001110110" => data <= triangle_rom(3702);
     when "111001110111" => data <= triangle_rom(3703);
     when "111001111000" => data <= triangle_rom(3704);
     when "111001111001" => data <= triangle_rom(3705);
     when "111001111010" => data <= triangle_rom(3706);
     when "111001111011" => data <= triangle_rom(3707);
     when "111001111100" => data <= triangle_rom(3708);
     when "111001111101" => data <= triangle_rom(3709);
     when "111001111110" => data <= triangle_rom(3710);
     when "111001111111" => data <= triangle_rom(3711);
     when "111010000000" => data <= triangle_rom(3712);
     when "111010000001" => data <= triangle_rom(3713);
     when "111010000010" => data <= triangle_rom(3714);
     when "111010000011" => data <= triangle_rom(3715);
     when "111010000100" => data <= triangle_rom(3716);
     when "111010000101" => data <= triangle_rom(3717);
     when "111010000110" => data <= triangle_rom(3718);
     when "111010000111" => data <= triangle_rom(3719);
     when "111010001000" => data <= triangle_rom(3720);
     when "111010001001" => data <= triangle_rom(3721);
     when "111010001010" => data <= triangle_rom(3722);
     when "111010001011" => data <= triangle_rom(3723);
     when "111010001100" => data <= triangle_rom(3724);
     when "111010001101" => data <= triangle_rom(3725);
     when "111010001110" => data <= triangle_rom(3726);
     when "111010001111" => data <= triangle_rom(3727);
     when "111010010000" => data <= triangle_rom(3728);
     when "111010010001" => data <= triangle_rom(3729);
     when "111010010010" => data <= triangle_rom(3730);
     when "111010010011" => data <= triangle_rom(3731);
     when "111010010100" => data <= triangle_rom(3732);
     when "111010010101" => data <= triangle_rom(3733);
     when "111010010110" => data <= triangle_rom(3734);
     when "111010010111" => data <= triangle_rom(3735);
     when "111010011000" => data <= triangle_rom(3736);
     when "111010011001" => data <= triangle_rom(3737);
     when "111010011010" => data <= triangle_rom(3738);
     when "111010011011" => data <= triangle_rom(3739);
     when "111010011100" => data <= triangle_rom(3740);
     when "111010011101" => data <= triangle_rom(3741);
     when "111010011110" => data <= triangle_rom(3742);
     when "111010011111" => data <= triangle_rom(3743);
     when "111010100000" => data <= triangle_rom(3744);
     when "111010100001" => data <= triangle_rom(3745);
     when "111010100010" => data <= triangle_rom(3746);
     when "111010100011" => data <= triangle_rom(3747);
     when "111010100100" => data <= triangle_rom(3748);
     when "111010100101" => data <= triangle_rom(3749);
     when "111010100110" => data <= triangle_rom(3750);
     when "111010100111" => data <= triangle_rom(3751);
     when "111010101000" => data <= triangle_rom(3752);
     when "111010101001" => data <= triangle_rom(3753);
     when "111010101010" => data <= triangle_rom(3754);
     when "111010101011" => data <= triangle_rom(3755);
     when "111010101100" => data <= triangle_rom(3756);
     when "111010101101" => data <= triangle_rom(3757);
     when "111010101110" => data <= triangle_rom(3758);
     when "111010101111" => data <= triangle_rom(3759);
     when "111010110000" => data <= triangle_rom(3760);
     when "111010110001" => data <= triangle_rom(3761);
     when "111010110010" => data <= triangle_rom(3762);
     when "111010110011" => data <= triangle_rom(3763);
     when "111010110100" => data <= triangle_rom(3764);
     when "111010110101" => data <= triangle_rom(3765);
     when "111010110110" => data <= triangle_rom(3766);
     when "111010110111" => data <= triangle_rom(3767);
     when "111010111000" => data <= triangle_rom(3768);
     when "111010111001" => data <= triangle_rom(3769);
     when "111010111010" => data <= triangle_rom(3770);
     when "111010111011" => data <= triangle_rom(3771);
     when "111010111100" => data <= triangle_rom(3772);
     when "111010111101" => data <= triangle_rom(3773);
     when "111010111110" => data <= triangle_rom(3774);
     when "111010111111" => data <= triangle_rom(3775);
     when "111011000000" => data <= triangle_rom(3776);
     when "111011000001" => data <= triangle_rom(3777);
     when "111011000010" => data <= triangle_rom(3778);
     when "111011000011" => data <= triangle_rom(3779);
     when "111011000100" => data <= triangle_rom(3780);
     when "111011000101" => data <= triangle_rom(3781);
     when "111011000110" => data <= triangle_rom(3782);
     when "111011000111" => data <= triangle_rom(3783);
     when "111011001000" => data <= triangle_rom(3784);
     when "111011001001" => data <= triangle_rom(3785);
     when "111011001010" => data <= triangle_rom(3786);
     when "111011001011" => data <= triangle_rom(3787);
     when "111011001100" => data <= triangle_rom(3788);
     when "111011001101" => data <= triangle_rom(3789);
     when "111011001110" => data <= triangle_rom(3790);
     when "111011001111" => data <= triangle_rom(3791);
     when "111011010000" => data <= triangle_rom(3792);
     when "111011010001" => data <= triangle_rom(3793);
     when "111011010010" => data <= triangle_rom(3794);
     when "111011010011" => data <= triangle_rom(3795);
     when "111011010100" => data <= triangle_rom(3796);
     when "111011010101" => data <= triangle_rom(3797);
     when "111011010110" => data <= triangle_rom(3798);
     when "111011010111" => data <= triangle_rom(3799);
     when "111011011000" => data <= triangle_rom(3800);
     when "111011011001" => data <= triangle_rom(3801);
     when "111011011010" => data <= triangle_rom(3802);
     when "111011011011" => data <= triangle_rom(3803);
     when "111011011100" => data <= triangle_rom(3804);
     when "111011011101" => data <= triangle_rom(3805);
     when "111011011110" => data <= triangle_rom(3806);
     when "111011011111" => data <= triangle_rom(3807);
     when "111011100000" => data <= triangle_rom(3808);
     when "111011100001" => data <= triangle_rom(3809);
     when "111011100010" => data <= triangle_rom(3810);
     when "111011100011" => data <= triangle_rom(3811);
     when "111011100100" => data <= triangle_rom(3812);
     when "111011100101" => data <= triangle_rom(3813);
     when "111011100110" => data <= triangle_rom(3814);
     when "111011100111" => data <= triangle_rom(3815);
     when "111011101000" => data <= triangle_rom(3816);
     when "111011101001" => data <= triangle_rom(3817);
     when "111011101010" => data <= triangle_rom(3818);
     when "111011101011" => data <= triangle_rom(3819);
     when "111011101100" => data <= triangle_rom(3820);
     when "111011101101" => data <= triangle_rom(3821);
     when "111011101110" => data <= triangle_rom(3822);
     when "111011101111" => data <= triangle_rom(3823);
     when "111011110000" => data <= triangle_rom(3824);
     when "111011110001" => data <= triangle_rom(3825);
     when "111011110010" => data <= triangle_rom(3826);
     when "111011110011" => data <= triangle_rom(3827);
     when "111011110100" => data <= triangle_rom(3828);
     when "111011110101" => data <= triangle_rom(3829);
     when "111011110110" => data <= triangle_rom(3830);
     when "111011110111" => data <= triangle_rom(3831);
     when "111011111000" => data <= triangle_rom(3832);
     when "111011111001" => data <= triangle_rom(3833);
     when "111011111010" => data <= triangle_rom(3834);
     when "111011111011" => data <= triangle_rom(3835);
     when "111011111100" => data <= triangle_rom(3836);
     when "111011111101" => data <= triangle_rom(3837);
     when "111011111110" => data <= triangle_rom(3838);
     when "111011111111" => data <= triangle_rom(3839);
     when "111100000000" => data <= triangle_rom(3840);
     when "111100000001" => data <= triangle_rom(3841);
     when "111100000010" => data <= triangle_rom(3842);
     when "111100000011" => data <= triangle_rom(3843);
     when "111100000100" => data <= triangle_rom(3844);
     when "111100000101" => data <= triangle_rom(3845);
     when "111100000110" => data <= triangle_rom(3846);
     when "111100000111" => data <= triangle_rom(3847);
     when "111100001000" => data <= triangle_rom(3848);
     when "111100001001" => data <= triangle_rom(3849);
     when "111100001010" => data <= triangle_rom(3850);
     when "111100001011" => data <= triangle_rom(3851);
     when "111100001100" => data <= triangle_rom(3852);
     when "111100001101" => data <= triangle_rom(3853);
     when "111100001110" => data <= triangle_rom(3854);
     when "111100001111" => data <= triangle_rom(3855);
     when "111100010000" => data <= triangle_rom(3856);
     when "111100010001" => data <= triangle_rom(3857);
     when "111100010010" => data <= triangle_rom(3858);
     when "111100010011" => data <= triangle_rom(3859);
     when "111100010100" => data <= triangle_rom(3860);
     when "111100010101" => data <= triangle_rom(3861);
     when "111100010110" => data <= triangle_rom(3862);
     when "111100010111" => data <= triangle_rom(3863);
     when "111100011000" => data <= triangle_rom(3864);
     when "111100011001" => data <= triangle_rom(3865);
     when "111100011010" => data <= triangle_rom(3866);
     when "111100011011" => data <= triangle_rom(3867);
     when "111100011100" => data <= triangle_rom(3868);
     when "111100011101" => data <= triangle_rom(3869);
     when "111100011110" => data <= triangle_rom(3870);
     when "111100011111" => data <= triangle_rom(3871);
     when "111100100000" => data <= triangle_rom(3872);
     when "111100100001" => data <= triangle_rom(3873);
     when "111100100010" => data <= triangle_rom(3874);
     when "111100100011" => data <= triangle_rom(3875);
     when "111100100100" => data <= triangle_rom(3876);
     when "111100100101" => data <= triangle_rom(3877);
     when "111100100110" => data <= triangle_rom(3878);
     when "111100100111" => data <= triangle_rom(3879);
     when "111100101000" => data <= triangle_rom(3880);
     when "111100101001" => data <= triangle_rom(3881);
     when "111100101010" => data <= triangle_rom(3882);
     when "111100101011" => data <= triangle_rom(3883);
     when "111100101100" => data <= triangle_rom(3884);
     when "111100101101" => data <= triangle_rom(3885);
     when "111100101110" => data <= triangle_rom(3886);
     when "111100101111" => data <= triangle_rom(3887);
     when "111100110000" => data <= triangle_rom(3888);
     when "111100110001" => data <= triangle_rom(3889);
     when "111100110010" => data <= triangle_rom(3890);
     when "111100110011" => data <= triangle_rom(3891);
     when "111100110100" => data <= triangle_rom(3892);
     when "111100110101" => data <= triangle_rom(3893);
     when "111100110110" => data <= triangle_rom(3894);
     when "111100110111" => data <= triangle_rom(3895);
     when "111100111000" => data <= triangle_rom(3896);
     when "111100111001" => data <= triangle_rom(3897);
     when "111100111010" => data <= triangle_rom(3898);
     when "111100111011" => data <= triangle_rom(3899);
     when "111100111100" => data <= triangle_rom(3900);
     when "111100111101" => data <= triangle_rom(3901);
     when "111100111110" => data <= triangle_rom(3902);
     when "111100111111" => data <= triangle_rom(3903);
     when "111101000000" => data <= triangle_rom(3904);
     when "111101000001" => data <= triangle_rom(3905);
     when "111101000010" => data <= triangle_rom(3906);
     when "111101000011" => data <= triangle_rom(3907);
     when "111101000100" => data <= triangle_rom(3908);
     when "111101000101" => data <= triangle_rom(3909);
     when "111101000110" => data <= triangle_rom(3910);
     when "111101000111" => data <= triangle_rom(3911);
     when "111101001000" => data <= triangle_rom(3912);
     when "111101001001" => data <= triangle_rom(3913);
     when "111101001010" => data <= triangle_rom(3914);
     when "111101001011" => data <= triangle_rom(3915);
     when "111101001100" => data <= triangle_rom(3916);
     when "111101001101" => data <= triangle_rom(3917);
     when "111101001110" => data <= triangle_rom(3918);
     when "111101001111" => data <= triangle_rom(3919);
     when "111101010000" => data <= triangle_rom(3920);
     when "111101010001" => data <= triangle_rom(3921);
     when "111101010010" => data <= triangle_rom(3922);
     when "111101010011" => data <= triangle_rom(3923);
     when "111101010100" => data <= triangle_rom(3924);
     when "111101010101" => data <= triangle_rom(3925);
     when "111101010110" => data <= triangle_rom(3926);
     when "111101010111" => data <= triangle_rom(3927);
     when "111101011000" => data <= triangle_rom(3928);
     when "111101011001" => data <= triangle_rom(3929);
     when "111101011010" => data <= triangle_rom(3930);
     when "111101011011" => data <= triangle_rom(3931);
     when "111101011100" => data <= triangle_rom(3932);
     when "111101011101" => data <= triangle_rom(3933);
     when "111101011110" => data <= triangle_rom(3934);
     when "111101011111" => data <= triangle_rom(3935);
     when "111101100000" => data <= triangle_rom(3936);
     when "111101100001" => data <= triangle_rom(3937);
     when "111101100010" => data <= triangle_rom(3938);
     when "111101100011" => data <= triangle_rom(3939);
     when "111101100100" => data <= triangle_rom(3940);
     when "111101100101" => data <= triangle_rom(3941);
     when "111101100110" => data <= triangle_rom(3942);
     when "111101100111" => data <= triangle_rom(3943);
     when "111101101000" => data <= triangle_rom(3944);
     when "111101101001" => data <= triangle_rom(3945);
     when "111101101010" => data <= triangle_rom(3946);
     when "111101101011" => data <= triangle_rom(3947);
     when "111101101100" => data <= triangle_rom(3948);
     when "111101101101" => data <= triangle_rom(3949);
     when "111101101110" => data <= triangle_rom(3950);
     when "111101101111" => data <= triangle_rom(3951);
     when "111101110000" => data <= triangle_rom(3952);
     when "111101110001" => data <= triangle_rom(3953);
     when "111101110010" => data <= triangle_rom(3954);
     when "111101110011" => data <= triangle_rom(3955);
     when "111101110100" => data <= triangle_rom(3956);
     when "111101110101" => data <= triangle_rom(3957);
     when "111101110110" => data <= triangle_rom(3958);
     when "111101110111" => data <= triangle_rom(3959);
     when "111101111000" => data <= triangle_rom(3960);
     when "111101111001" => data <= triangle_rom(3961);
     when "111101111010" => data <= triangle_rom(3962);
     when "111101111011" => data <= triangle_rom(3963);
     when "111101111100" => data <= triangle_rom(3964);
     when "111101111101" => data <= triangle_rom(3965);
     when "111101111110" => data <= triangle_rom(3966);
     when "111101111111" => data <= triangle_rom(3967);
     when "111110000000" => data <= triangle_rom(3968);
     when "111110000001" => data <= triangle_rom(3969);
     when "111110000010" => data <= triangle_rom(3970);
     when "111110000011" => data <= triangle_rom(3971);
     when "111110000100" => data <= triangle_rom(3972);
     when "111110000101" => data <= triangle_rom(3973);
     when "111110000110" => data <= triangle_rom(3974);
     when "111110000111" => data <= triangle_rom(3975);
     when "111110001000" => data <= triangle_rom(3976);
     when "111110001001" => data <= triangle_rom(3977);
     when "111110001010" => data <= triangle_rom(3978);
     when "111110001011" => data <= triangle_rom(3979);
     when "111110001100" => data <= triangle_rom(3980);
     when "111110001101" => data <= triangle_rom(3981);
     when "111110001110" => data <= triangle_rom(3982);
     when "111110001111" => data <= triangle_rom(3983);
     when "111110010000" => data <= triangle_rom(3984);
     when "111110010001" => data <= triangle_rom(3985);
     when "111110010010" => data <= triangle_rom(3986);
     when "111110010011" => data <= triangle_rom(3987);
     when "111110010100" => data <= triangle_rom(3988);
     when "111110010101" => data <= triangle_rom(3989);
     when "111110010110" => data <= triangle_rom(3990);
     when "111110010111" => data <= triangle_rom(3991);
     when "111110011000" => data <= triangle_rom(3992);
     when "111110011001" => data <= triangle_rom(3993);
     when "111110011010" => data <= triangle_rom(3994);
     when "111110011011" => data <= triangle_rom(3995);
     when "111110011100" => data <= triangle_rom(3996);
     when "111110011101" => data <= triangle_rom(3997);
     when "111110011110" => data <= triangle_rom(3998);
     when "111110011111" => data <= triangle_rom(3999);
     when "111110100000" => data <= triangle_rom(4000);
     when "111110100001" => data <= triangle_rom(4001);
     when "111110100010" => data <= triangle_rom(4002);
     when "111110100011" => data <= triangle_rom(4003);
     when "111110100100" => data <= triangle_rom(4004);
     when "111110100101" => data <= triangle_rom(4005);
     when "111110100110" => data <= triangle_rom(4006);
     when "111110100111" => data <= triangle_rom(4007);
     when "111110101000" => data <= triangle_rom(4008);
     when "111110101001" => data <= triangle_rom(4009);
     when "111110101010" => data <= triangle_rom(4010);
     when "111110101011" => data <= triangle_rom(4011);
     when "111110101100" => data <= triangle_rom(4012);
     when "111110101101" => data <= triangle_rom(4013);
     when "111110101110" => data <= triangle_rom(4014);
     when "111110101111" => data <= triangle_rom(4015);
     when "111110110000" => data <= triangle_rom(4016);
     when "111110110001" => data <= triangle_rom(4017);
     when "111110110010" => data <= triangle_rom(4018);
     when "111110110011" => data <= triangle_rom(4019);
     when "111110110100" => data <= triangle_rom(4020);
     when "111110110101" => data <= triangle_rom(4021);
     when "111110110110" => data <= triangle_rom(4022);
     when "111110110111" => data <= triangle_rom(4023);
     when "111110111000" => data <= triangle_rom(4024);
     when "111110111001" => data <= triangle_rom(4025);
     when "111110111010" => data <= triangle_rom(4026);
     when "111110111011" => data <= triangle_rom(4027);
     when "111110111100" => data <= triangle_rom(4028);
     when "111110111101" => data <= triangle_rom(4029);
     when "111110111110" => data <= triangle_rom(4030);
     when "111110111111" => data <= triangle_rom(4031);
     when "111111000000" => data <= triangle_rom(4032);
     when "111111000001" => data <= triangle_rom(4033);
     when "111111000010" => data <= triangle_rom(4034);
     when "111111000011" => data <= triangle_rom(4035);
     when "111111000100" => data <= triangle_rom(4036);
     when "111111000101" => data <= triangle_rom(4037);
     when "111111000110" => data <= triangle_rom(4038);
     when "111111000111" => data <= triangle_rom(4039);
     when "111111001000" => data <= triangle_rom(4040);
     when "111111001001" => data <= triangle_rom(4041);
     when "111111001010" => data <= triangle_rom(4042);
     when "111111001011" => data <= triangle_rom(4043);
     when "111111001100" => data <= triangle_rom(4044);
     when "111111001101" => data <= triangle_rom(4045);
     when "111111001110" => data <= triangle_rom(4046);
     when "111111001111" => data <= triangle_rom(4047);
     when "111111010000" => data <= triangle_rom(4048);
     when "111111010001" => data <= triangle_rom(4049);
     when "111111010010" => data <= triangle_rom(4050);
     when "111111010011" => data <= triangle_rom(4051);
     when "111111010100" => data <= triangle_rom(4052);
     when "111111010101" => data <= triangle_rom(4053);
     when "111111010110" => data <= triangle_rom(4054);
     when "111111010111" => data <= triangle_rom(4055);
     when "111111011000" => data <= triangle_rom(4056);
     when "111111011001" => data <= triangle_rom(4057);
     when "111111011010" => data <= triangle_rom(4058);
     when "111111011011" => data <= triangle_rom(4059);
     when "111111011100" => data <= triangle_rom(4060);
     when "111111011101" => data <= triangle_rom(4061);
     when "111111011110" => data <= triangle_rom(4062);
     when "111111011111" => data <= triangle_rom(4063);
     when "111111100000" => data <= triangle_rom(4064);
     when "111111100001" => data <= triangle_rom(4065);
     when "111111100010" => data <= triangle_rom(4066);
     when "111111100011" => data <= triangle_rom(4067);
     when "111111100100" => data <= triangle_rom(4068);
     when "111111100101" => data <= triangle_rom(4069);
     when "111111100110" => data <= triangle_rom(4070);
     when "111111100111" => data <= triangle_rom(4071);
     when "111111101000" => data <= triangle_rom(4072);
     when "111111101001" => data <= triangle_rom(4073);
     when "111111101010" => data <= triangle_rom(4074);
     when "111111101011" => data <= triangle_rom(4075);
     when "111111101100" => data <= triangle_rom(4076);
     when "111111101101" => data <= triangle_rom(4077);
     when "111111101110" => data <= triangle_rom(4078);
     when "111111101111" => data <= triangle_rom(4079);
     when "111111110000" => data <= triangle_rom(4080);
     when "111111110001" => data <= triangle_rom(4081);
     when "111111110010" => data <= triangle_rom(4082);
     when "111111110011" => data <= triangle_rom(4083);
     when "111111110100" => data <= triangle_rom(4084);
     when "111111110101" => data <= triangle_rom(4085);
     when "111111110110" => data <= triangle_rom(4086);
     when "111111110111" => data <= triangle_rom(4087);
     when "111111111000" => data <= triangle_rom(4088);
     when "111111111001" => data <= triangle_rom(4089);
     when "111111111010" => data <= triangle_rom(4090);
     when "111111111011" => data <= triangle_rom(4091);
     when "111111111100" => data <= triangle_rom(4092);
     when "111111111101" => data <= triangle_rom(4093);
     when "111111111110" => data <= triangle_rom(4094);
     when "111111111111" => data <= triangle_rom(4095);
     when others => data <= "000000000000";
    end case;
 end process;
end arch_Triangle_LUT;
